`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    12:13:19 09/20/2021 
// Design Name: 
// Module Name:    RL_Int 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module RL_Int(
	input clk, rst,
	input signed [31:0] Signal,
	output reg signed [31:0] Output,
	output reg OutInd
    );
    parameter Wind = 32;
integer f1;
reg signed [31:0] Reg [0:Wind-1];
reg signed [63:0]  sum;
reg signed [31:0]  temp;
reg signed [63:0] temp1;
reg signed[31:0] Coff [0:Wind-1];

integer i =0;


initial begin

for (i=0; i<Wind;i=i+1)
begin
	Reg[i] =0;
end
OutInd = 0;

//Coff[127]=83828.3083224284;
//Coff[126]=84158.9958363417;
//Coff[125]=84493.6280104285;
//Coff[124]=84832.2838981899;
//Coff[123]=85175.0447890604;
//Coff[122]=85521.9942904109;
//Coff[121]=85873.2184131728;
//Coff[120]=86228.8056614541;
//Coff[119]=86588.8471262248;
//Coff[118]=86953.4365833365;
//Coff[117]=87322.6705961562;
//Coff[116]=87696.648623002;
//Coff[115]=88075.4731296767;
//Coff[114]=88459.2497074565;
//Coff[113]=88848.0871967083;
//Coff[112]=89242.0978165845;
//Coff[111]=89641.3973010861;
//Coff[110]=90046.1050418824;
//Coff[109]=90456.3442383101;
//Coff[108]=90872.2420549186;
//Coff[107]=91293.9297870862;
//Coff[106]=91721.5430351775;
//Coff[105]=92155.221887724;
//Coff[104]=92595.1111142587;
//Coff[103]=93041.3603683606;
//Coff[102]=93494.1244015644;
//Coff[101]=93953.5632888319;
//Coff[100]=94419.8426663509;
//Coff[99]=94893.1339824262;
//Coff[98]=95373.6147623532;
//Coff[97]=95861.4688882053;
//Coff[96]=96356.8868945044;
//Coff[95]=96860.0662809101;
//Coff[94]=97371.2118430252;
//Coff[93]=97890.5360226482;
//Coff[92]=98418.2592787434;
//Coff[91]=98954.6104807182;
//Coff[90]=99499.8273254947;
//Coff[89]=100054.156780142;
//Coff[88]=100617.855551951;
//Coff[87]=101191.190588001;
//Coff[86]=101774.439606344;
//Coff[85]=102367.891661318;
//Coff[84]=102971.847745526;
//Coff[83]=103586.621431353;
//Coff[82]=104212.539555135;
//Coff[81]=104849.942947352;
//Coff[80]=105499.187212563;
//Coff[79]=106160.643563163;
//Coff[78]=106834.699711323;
//Coff[77]=107521.760824102;
//Coff[76]=108222.250546941;
//Coff[75]=108936.612101546;
//Coff[74]=109665.309464516;
//Coff[73]=110408.828633902;
//Coff[72]=111167.678991536;
//Coff[71]=111942.394769794;
//Coff[70]=112733.536632415;
//Coff[69]=113541.693379962;
//Coff[68]=114367.483791792;
//Coff[67]=115211.55861754;
//Coff[66]=116074.602732745;
//Coff[65]=116957.337474822;
//Coff[64]=117860.523177488;
//Coff[63]=118784.961923912;
//Coff[62]=119731.500541179;
//Coff[61]=120701.033861562;
//Coff[60]=121694.508279097;
//Coff[59]=122712.925633631;
//Coff[58]=123757.347458518;
//Coff[57]=124828.899633026;
//Coff[56]=125928.777485667;
//Coff[55]=127058.251401186;
//Coff[54]=128218.672990912;
//Coff[53]=129411.481894686;
//Coff[52]=130638.213292173;
//Coff[51]=131900.506212733;
//Coff[50]=133200.112746117;
//Coff[49]=134538.908271751;
//Coff[48]=135918.902842482;
//Coff[47]=137342.253879967;
//Coff[46]=138811.280364173;
//Coff[45]=140328.478729338;
//Coff[44]=141896.540714374;
//Coff[43]=143518.373458222;
//Coff[42]=145197.122181657;
//Coff[41]=146936.195858423;
//Coff[40]=148739.296352766;
//Coff[39]=150610.451590547;
//Coff[38]=152554.053440853;
//Coff[37]=154574.90111977;
//Coff[36]=156678.251093578;
//Coff[35]=158869.874663907;
//Coff[34]=161156.124672794;
//Coff[33]=163544.013085393;
//Coff[32]=166041.301610965;
Coff[31]=168656.608033694;
Coff[30]=171399.531577049;
Coff[29]=174280.80146436;
Coff[28]=177312.453925213;
Coff[27]=180508.044318099;
Coff[26]=183882.902912123;
Coff[25]=187454.445362554;
Coff[24]=191242.552263745;
Coff[23]=195270.036712663;
Coff[22]=199563.225069153;
Coff[21]=204152.684800594;
Coff[20]=209074.145573202;
Coff[19]=214369.677322765;
Coff[18]=220089.21459575;
Coff[17]=226292.554286982;
Coff[16]=233052.011001298;
Coff[15]=240456.002302875;
Coff[14]=248613.975105421;
Coff[13]=257663.309789479;
Coff[12]=267779.215036541;
Coff[11]=279189.276843926;
Coff[10]=292195.493925534;
Coff[9]=307208.828622374;
Coff[8]=324805.65701653;
Coff[7]=345824.697500158;
Coff[6]=371543.97242826;
Coff[5]=404030.046077806;
Coff[4]=446901.728603397;
Coff[3]=507256.251117158;
Coff[2]=601699.628204182;
Coff[1]=784150.222304811;
Coff[0]=1893106.10162615;

	f1 = $fopen("Output.txt") ;

end

always @(posedge clk)
begin
	if (rst ==0)
	begin
	
		for (i=1; i<Wind; i=i+1)
		begin
			Reg[i-1] = Reg[i];
			$monitor("Reg[%d]= %d \n" , i,$signed(Reg[i]) ) ;
		end
		// New Input at last position (31)
		Reg[Wind-1]= Signal;
		$monitor("Reg[%d]= %d \n" , i,$signed(Reg[i]) ) ;
		
		sum =0;
		// Add every two adjasent signals to each other and average them 
		for (i=0; i<Wind-1; i=i+1)
		begin
		// reg[31]  
			temp = (Reg[i+1] + Reg[i]);
//			$monitor("temp= %d \n" ,$signed(temp) ) ;
			temp = temp >>> 1;
//			$monitor("coff= %d \n" ,$signed(Coff[Wind-1-i]) ) ;
			temp1 = temp * Coff[Wind-1-i];
			sum = sum + temp1[55:24];
			$monitor("sum= %d \n" ,$signed(sum) ) ;
		end
		Output = sum[31:0];
		OutInd = !OutInd;
		
		
	end

end

endmodule
