

module IIR_PhasOpti(

input clk, rst,
input signed [31:0] Signal,
output reg signed [31:0] Output,
output reg OutInd
);

parameter N = 8;

  reg signed [31:0] aCoff[0:N];
    reg signed [31:0] bCoff[0:N];
    reg signed [31:0] RegA[0:N-1];
     reg signed [31:0] RegB[0:N-1];
     reg signed [64:0] sum;
     reg signed [63:0]temp ;
     reg signed [31:0]temp1 ;
     reg signed [96:0]temp2;
     reg signed [31:0] MagDiff;
integer i =0;
integer j =0;
integer k =0;

    
  
//reg signed [63:0] temp;
//reg signed [31:0] temp1;
//reg signed [31:0] temp2;
//reg signed [31:0] PrevSig;
//integer StepBeta = 16861102;
//integer alpha = 8388608; // .5 *2^24
//integer step =   167770; // .01 *2^24
//integer beta = 8388608; // (1- alpha)


initial 
begin
//PrevSig = 0;
//OutInd = 0;



        // 5th Order IIR //////////////////////////////////////////////////////
        /////////////////////////////////////////////////////////////////////////
        //    MagDiff = 342171;
//        aCoff[0] = 16777216;
//        aCoff[1] = 78901;
//        aCoff[2] = -5612413;
//        aCoff[3] = 1932272;
//        aCoff[4] = -7936566;
//        aCoff[5] = -1610345;
        
//        bCoff[0] = 14579422;
//        bCoff[1] = 14579422;
//        bCoff[2] = 2318216;
//        bCoff[3] = 4326682;
//        bCoff[4] = -1711277;
//        bCoff[5] = -3807764;
////////////////////////////////////////////


        // 3r Order IIR //////////////////////////////////////////////////////
        /////////////////////////////////////////////////////////////////////////
//            MagDiff = 3562675.37269376;
//     bCoff[0] =8877736.68384249;
//     bCoff[1] =	2437411.98466256;
//  	 bCoff[2] =-7136437.70922856;
//  	 bCoff[3]=	-1268239.59577874;
  	 
////  	 bCoff[4] =-6239235.70922856;
////        bCoff[5]=    2430269.59577874;
  	 
  				
//    aCoff[0] =16777216;
//    aCoff[1] =    -12192520.4347745;
//    aCoff[2] =-9972937.18397900;
//    aCoff[3]=    5697900.32590527 ;
    
    
    
    ////////////////////////////////
    
    // 5th order derivtive
    
//     MagDiff = 3562675.37269376;
//    bCoff[0] =16777216;
//      bCoff[1] =	-10258798.6752615;
//      bCoff[2] =	6108101.45446478; 
//      bCoff[3] =	-3725243.39955478	;
//      bCoff[4] =-10778461.4688899; 
//      bCoff[5] =	3456125.69763234;
      
//        aCoff[0] =16777216 ;  
//     aCoff[1] =6504047.96376353 ;  
//     aCoff[2] = 4266704.69527860 ;  
//     aCoff[3] = 5551333.39800030;
//     aCoff[4] =    -10359961.9354427 ;
//     aCoff[5] =   -3193439.81394206;
     
     
     /////////////////////////////////
//     5th order integral
//16777216	14547578.9957828	12383937.0244806	14761680.6362237	-323272.578163656	-2121234.29765006
//16777216	-2649206.52514009	5528668.05103169	194773.218047348	-9948210.92583126	-1866144.18311735

//MagDiff = 3562675.37269376;
//      bCoff[0] =16777216;
//     bCoff[1] =   14547578.9957828;
//     bCoff[2] =   12383937.0244806; 
//     bCoff[3] =   14761680.6362237    ;
//     bCoff[4] =-323272.578163656; 
//     bCoff[5] =   -2121234.29765006;
     
//       aCoff[0] =16777216 ;  
//    aCoff[1] = -2649206.52514009 ;  
//    aCoff[2] = 5528668.05103169 ;  
//    aCoff[3] =  194773.218047348;
//    aCoff[4] = -9948210.92583126;
//     aCoff[5] =   -1866144.18311735;
////     aCoff[4] =    -1116752.4347745;
//       aCoff[5] =-567293.18397900;
//       aCoff[3]=    5697900.32590527 ;
    
//       3r Order IIR Diff .5 //////////////////////////////////////////////////////
          /////////////////////////////////////////////////////////////////////
//         MagDiff =  156052427;
  
//       bCoff[0] =16777216;
//       bCoff[1] =   -9607942.80347991;
//         bCoff[2] =-11558591.3889144;
//         bCoff[3]=    4871167.15444841;
         
                    
//      aCoff[0] =16777216;
//      aCoff[1] =   7251861.71295358;
//      aCoff[2] =-12637330.0249737;
//      aCoff[3]=   -3822578.32928449 ;


////////// 3rd derivative

//  MagDiff =  156052427;
  
//       bCoff[0] =16777216;
//       bCoff[1] =  13806676.9425647 ;
//         bCoff[2] =  -8822890.85827767  ;
//         bCoff[3]=    -6084491.85362399;
         
                    
//      aCoff[0] =16777216;
//      aCoff[1] =   -2974507.69031855  ;
//      aCoff[2] =-13871752.8172013;
//      aCoff[3]=   1460634.19887561 ;

// //////////////////////////////////////////////////////////
///////////////////////////////////////////////////////////   8th order integral
MagDiff =  156052427;
bCoff[0] =16777216 ;
bCoff[1] =	14926961.6327024  ;
bCoff[2] =	-6357951.88273083  ;
bCoff[3] =	-11437820.6255520 ;
bCoff[4] =	-9939972.91105323 ;
bCoff[5] =	-6030294.75185011 ;
bCoff[6] =	-5267598.64578749	 ;
bCoff[7] =3223333.14044006	 ;
bCoff[8] =5487085.29799556;
 
 aCoff[0] =16777216	;
  aCoff[1] = -823710.280681265	; 
  aCoff[2] = -13319594.0772525	; 
  aCoff[3] = -7294901.82814357;
   aCoff[4] = 	-1869618.06647181; 
   aCoff[5] = 	1558566.48948471	;
    aCoff[6] = -2730698.52227539; 
    aCoff[7] = 	5908846.12869325;
     aCoff[8] = 	1874996.36923806;
     
     // //////////////////////////////////////////////////////////
     ///////////////////////////////////////////////////////////   8th order Derivative
     MagDiff =  156052427;
     bCoff[0] =16777216 ;
     bCoff[1] =   -4624124.60436625;
     bCoff[2] =   2012996.26737830  ;
     bCoff[3] =    -5842851.46645201 ;
     bCoff[4] =   -4636056.01738069;
     bCoff[5] =   1510867.30008868 ;
     bCoff[6] =    -664136.274307931    ;
     bCoff[7] =-164698.238328802     ;
     bCoff[8] =-1649678.0726699;
      
      aCoff[0] =16777216    ;
       aCoff[1] = 12094566.5926713      ; 
       aCoff[2] = 5755406.03237154     ; 
       aCoff[3] = 2298439.32473590;
        aCoff[4] =    -5391104.52342875; 
        aCoff[5] =    -404491.197662144    ;
         aCoff[6] = 8479.64832957476; 
         aCoff[7] =     557308.287966320;
          aCoff[8] =    -1000080.14499001;
        for(i = 0; i<=N-1; i= i+1) begin
            RegA[i] =0;
            RegB[i] = 0;
        end
        

        
        
end
always @ (posedge clk)
begin
    if (!rst)
    begin


           for (j = 0 ; j<=N ; j= j+1) begin
               if (j == 0) 
                 sum =   bCoff[j]*Signal;
               else
                 sum = sum+  bCoff[j]*RegB[j-1] ;     
               
           end
           
     

             for (j = N ; j>=0 ; j= j-1) begin
               if (j == 0) begin
               //    [96:0]  (25e72)    = (17e48)*(8e24);
                    temp2 = aCoff[j]*sum;
                    temp1 = temp2[79:48];
                     temp = temp1*MagDiff;
                    Output = temp[55:24];
                    if( Output == 135151) begin
                    Output = Output;
                    end
              end  else
                 sum = sum  - aCoff[j]*RegA[j-1];
                
             end
             
            for (k = N ; k>=0 ; k= k-1) begin
                        if (k == 0) begin
                          RegB[k] =   Signal;
                           RegA[k] =  temp1;
                       end  else
                        begin
                         RegB[k] = RegB[k-1] ;
                          RegA[k] = RegA[k-1] ;
                        end
                    end
    
       end
   
end

endmodule