`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    14:27:11 08/22/2021 
// Design Name: 
// Module Name:    SignalLUT 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module SignalLUT(

	input control,
   input  rst,
	output reg [31:0] Signal,
	output reg SigInd
    );
    
    parameter SigLength = 666;
	reg signed [31:0] Input [0:SigLength];
	 
	
	integer i=0;
	
initial begin



// Sin F =.15 Ts =.01
Input[	0	]=	0	;
Input[	1	]=	158119.1947	;
Input[	2	]=	316224.3444	;
Input[	3	]=	474301.4051	;
Input[	4	]=	632336.3357	;
Input[	5	]=	790315.0985	;
Input[	6	]=	948223.661	;
Input[	7	]=	1106047.997	;
Input[	8	]=	1263774.087	;
Input[	9	]=	1421387.921	;
Input[	10	]=	1578875.5	;
Input[	11	]=	1736222.834	;
Input[	12	]=	1893415.946	;
Input[	13	]=	2050440.874	;
Input[	14	]=	2207283.67	;
Input[	15	]=	2363930.403	;
Input[	16	]=	2520367.157	;
Input[	17	]=	2676580.038	;
Input[	18	]=	2832555.17	;
Input[	19	]=	2988278.698	;
Input[	20	]=	3143736.789	;
Input[	21	]=	3298915.636	;
Input[	22	]=	3453801.454	;
Input[	23	]=	3608380.485	;
Input[	24	]=	3762638.999	;
Input[	25	]=	3916563.294	;
Input[	26	]=	4070139.696	;
Input[	27	]=	4223354.566	;
Input[	28	]=	4376194.293	;
Input[	29	]=	4528645.301	;
Input[	30	]=	4680694.048	;
Input[	31	]=	4832327.029	;
Input[	32	]=	4983530.775	;
Input[	33	]=	5134291.855	;
Input[	34	]=	5284596.877	;
Input[	35	]=	5434432.491	;
Input[	36	]=	5583785.387	;
Input[	37	]=	5732642.3	;
Input[	38	]=	5880990.005	;
Input[	39	]=	6028815.327	;
Input[	40	]=	6176105.135	;
Input[	41	]=	6322846.346	;
Input[	42	]=	6469025.925	;
Input[	43	]=	6614630.887	;
Input[	44	]=	6759648.3	;
Input[	45	]=	6904065.281	;
Input[	46	]=	7047869.004	;
Input[	47	]=	7191046.694	;
Input[	48	]=	7333585.634	;
Input[	49	]=	7475473.162	;
Input[	50	]=	7616696.676	;
Input[	51	]=	7757243.631	;
Input[	52	]=	7897101.542	;
Input[	53	]=	8036257.987	;
Input[	54	]=	8174700.605	;
Input[	55	]=	8312417.099	;
Input[	56	]=	8449395.236	;
Input[	57	]=	8585622.849	;
Input[	58	]=	8721087.838	;
Input[	59	]=	8855778.169	;
Input[	60	]=	8989681.878	;
Input[	61	]=	9122787.072	;
Input[	62	]=	9255081.927	;
Input[	63	]=	9386554.692	;
Input[	64	]=	9517193.69	;
Input[	65	]=	9646987.315	;
Input[	66	]=	9775924.039	;
Input[	67	]=	9903992.408	;
Input[	68	]=	10031181.05	;
Input[	69	]=	10157478.66	;
Input[	70	]=	10282874.03	;
Input[	71	]=	10407356.01	;
Input[	72	]=	10530913.55	;
Input[	73	]=	10653535.67	;
Input[	74	]=	10775211.49	;
Input[	75	]=	10895930.19	;
Input[	76	]=	11015681.05	;
Input[	77	]=	11134453.43	;
Input[	78	]=	11252236.79	;
Input[	79	]=	11369020.65	;
Input[	80	]=	11484794.66	;
Input[	81	]=	11599548.52	;
Input[	82	]=	11713272.04	;
Input[	83	]=	11825955.12	;
Input[	84	]=	11937587.75	;
Input[	85	]=	12048160.01	;
Input[	86	]=	12157662.09	;
Input[	87	]=	12266084.25	;
Input[	88	]=	12373416.87	;
Input[	89	]=	12479650.41	;
Input[	90	]=	12584775.44	;
Input[	91	]=	12688782.61	;
Input[	92	]=	12791662.69	;
Input[	93	]=	12893406.55	;
Input[	94	]=	12994005.13	;
Input[	95	]=	13093449.52	;
Input[	96	]=	13191730.86	;
Input[	97	]=	13288840.45	;
Input[	98	]=	13384769.64	;
Input[	99	]=	13479509.91	;
Input[	100	]=	13573052.86	;
Input[	101	]=	13665390.17	;
Input[	102	]=	13756513.65	;
Input[	103	]=	13846415.19	;
Input[	104	]=	13935086.81	;
Input[	105	]=	14022520.64	;
Input[	106	]=	14108708.9	;
Input[	107	]=	14193643.95	;
Input[	108	]=	14277318.24	;
Input[	109	]=	14359724.33	;
Input[	110	]=	14440854.91	;
Input[	111	]=	14520702.77	;
Input[	112	]=	14599260.81	;
Input[	113	]=	14676522.07	;
Input[	114	]=	14752479.67	;
Input[	115	]=	14827126.87	;
Input[	116	]=	14900457.04	;
Input[	117	]=	14972463.66	;
Input[	118	]=	15043140.35	;
Input[	119	]=	15112480.81	;
Input[	120	]=	15180478.9	;
Input[	121	]=	15247128.57	;
Input[	122	]=	15312423.9	;
Input[	123	]=	15376359.1	;
Input[	124	]=	15438928.47	;
Input[	125	]=	15500126.47	;
Input[	126	]=	15559947.67	;
Input[	127	]=	15618386.73	;
Input[	128	]=	15675438.48	;
Input[	129	]=	15731097.85	;
Input[	130	]=	15785359.89	;
Input[	131	]=	15838219.78	;
Input[	132	]=	15889672.84	;
Input[	133	]=	15939714.47	;
Input[	134	]=	15988340.26	;
Input[	135	]=	16035545.86	;
Input[	136	]=	16081327.1	;
Input[	137	]=	16125679.89	;
Input[	138	]=	16168600.31	;
Input[	139	]=	16210084.55	;
Input[	140	]=	16250128.91	;
Input[	141	]=	16288729.84	;
Input[	142	]=	16325883.91	;
Input[	143	]=	16361587.82	;
Input[	144	]=	16395838.4	;
Input[	145	]=	16428632.61	;
Input[	146	]=	16459967.53	;
Input[	147	]=	16489840.38	;
Input[	148	]=	16518248.51	;
Input[	149	]=	16545189.39	;
Input[	150	]=	16570660.63	;
Input[	151	]=	16594659.97	;
Input[	152	]=	16617185.28	;
Input[	153	]=	16638234.55	;
Input[	154	]=	16657805.92	;
Input[	155	]=	16675897.65	;
Input[	156	]=	16692508.12	;
Input[	157	]=	16707635.87	;
Input[	158	]=	16721279.55	;
Input[	159	]=	16733437.96	;
Input[	160	]=	16744110	;
Input[	161	]=	16753294.73	;
Input[	162	]=	16760991.34	;
Input[	163	]=	16767199.14	;
Input[	164	]=	16771917.58	;
Input[	165	]=	16775146.24	;
Input[	166	]=	16776884.83	;
Input[	167	]=	16777133.21	;
Input[	168	]=	16775891.34	;
Input[	169	]=	16773159.34	;
Input[	170	]=	16768937.46	;
Input[	171	]=	16763226.06	;
Input[	172	]=	16756025.65	;
Input[	173	]=	16747336.87	;
Input[	174	]=	16737160.5	;
Input[	175	]=	16725497.44	;
Input[	176	]=	16712348.73	;
Input[	177	]=	16697715.52	;
Input[	178	]=	16681599.13	;
Input[	179	]=	16664000.98	;
Input[	180	]=	16644922.64	;
Input[	181	]=	16624365.8	;
Input[	182	]=	16602332.29	;
Input[	183	]=	16578824.06	;
Input[	184	]=	16553843.21	;
Input[	185	]=	16527391.95	;
Input[	186	]=	16499472.63	;
Input[	187	]=	16470087.73	;
Input[	188	]=	16439239.86	;
Input[	189	]=	16406931.77	;
Input[	190	]=	16373166.31	;
Input[	191	]=	16337946.5	;
Input[	192	]=	16301275.46	;
Input[	193	]=	16263156.44	;
Input[	194	]=	16223592.83	;
Input[	195	]=	16182588.15	;
Input[	196	]=	16140146.04	;
Input[	197	]=	16096270.27	;
Input[	198	]=	16050964.74	;
Input[	199	]=	16004233.46	;
Input[	200	]=	15956080.6	;
Input[	201	]=	15906510.43	;
Input[	202	]=	15855527.35	;
Input[	203	]=	15803135.88	;
Input[	204	]=	15749340.7	;
Input[	205	]=	15694146.56	;
Input[	206	]=	15637558.38	;
Input[	207	]=	15579581.18	;
Input[	208	]=	15520220.12	;
Input[	209	]=	15459480.45	;
Input[	210	]=	15397367.59	;
Input[	211	]=	15333887.04	;
Input[	212	]=	15269044.45	;
Input[	213	]=	15202845.58	;
Input[	214	]=	15135296.3	;
Input[	215	]=	15066402.61	;
Input[	216	]=	14996170.64	;
Input[	217	]=	14924606.63	;
Input[	218	]=	14851716.92	;
Input[	219	]=	14777508	;
Input[	220	]=	14701986.45	;
Input[	221	]=	14625158.99	;
Input[	222	]=	14547032.44	;
Input[	223	]=	14467613.74	;
Input[	224	]=	14386909.94	;
Input[	225	]=	14304928.21	;
Input[	226	]=	14221675.83	;
Input[	227	]=	14137160.21	;
Input[	228	]=	14051388.83	;
Input[	229	]=	13964369.34	;
Input[	230	]=	13876109.44	;
Input[	231	]=	13786616.99	;
Input[	232	]=	13695899.94	;
Input[	233	]=	13603966.33	;
Input[	234	]=	13510824.35	;
Input[	235	]=	13416482.25	;
Input[	236	]=	13320948.42	;
Input[	237	]=	13224231.35	;
Input[	238	]=	13126339.63	;
Input[	239	]=	13027281.94	;
Input[	240	]=	12927067.1	;
Input[	241	]=	12825704.01	;
Input[	242	]=	12723201.66	;
Input[	243	]=	12619569.16	;
Input[	244	]=	12514815.72	;
Input[	245	]=	12408950.64	;
Input[	246	]=	12301983.33	;
Input[	247	]=	12193923.28	;
Input[	248	]=	12084780.1	;
Input[	249	]=	11974563.48	;
Input[	250	]=	11863283.2	;
Input[	251	]=	11750949.17	;
Input[	252	]=	11637571.34	;
Input[	253	]=	11523159.8	;
Input[	254	]=	11407724.7	;
Input[	255	]=	11291276.31	;
Input[	256	]=	11173824.96	;
Input[	257	]=	11055381.08	;
Input[	258	]=	10935955.21	;
Input[	259	]=	10815557.93	;
Input[	260	]=	10694199.96	;
Input[	261	]=	10571892.07	;
Input[	262	]=	10448645.12	;
Input[	263	]=	10324470.06	;
Input[	264	]=	10199377.92	;
Input[	265	]=	10073379.81	;
Input[	266	]=	9946486.929	;
Input[	267	]=	9818710.542	;
Input[	268	]=	9690062.001	;
Input[	269	]=	9560552.732	;
Input[	270	]=	9430194.24	;
Input[	271	]=	9298998.104	;
Input[	272	]=	9166975.976	;
Input[	273	]=	9034139.585	;
Input[	274	]=	8900500.73	;
Input[	275	]=	8766071.28	;
Input[	276	]=	8630863.177	;
Input[	277	]=	8494888.431	;
Input[	278	]=	8358159.12	;
Input[	279	]=	8220687.389	;
Input[	280	]=	8082485.449	;
Input[	281	]=	7943565.576	;
Input[	282	]=	7803940.11	;
Input[	283	]=	7663621.452	;
Input[	284	]=	7522622.067	;
Input[	285	]=	7380954.48	;
Input[	286	]=	7238631.273	;
Input[	287	]=	7095665.089	;
Input[	288	]=	6952068.627	;
Input[	289	]=	6807854.643	;
Input[	290	]=	6663035.945	;
Input[	291	]=	6517625.398	;
Input[	292	]=	6371635.918	;
Input[	293	]=	6225080.472	;
Input[	294	]=	6077972.079	;
Input[	295	]=	5930323.805	;
Input[	296	]=	5782148.765	;
Input[	297	]=	5633460.121	;
Input[	298	]=	5484271.081	;
Input[	299	]=	5334594.897	;
Input[	300	]=	5184444.862	;
Input[	301	]=	5033834.316	;
Input[	302	]=	4882776.635	;
Input[	303	]=	4731285.237	;
Input[	304	]=	4579373.58	;
Input[	305	]=	4427055.156	;
Input[	306	]=	4274343.495	;
Input[	307	]=	4121252.163	;
Input[	308	]=	3967794.757	;
Input[	309	]=	3813984.908	;
Input[	310	]=	3659836.28	;
Input[	311	]=	3505362.563	;
Input[	312	]=	3350577.48	;
Input[	313	]=	3195494.78	;
Input[	314	]=	3040128.237	;
Input[	315	]=	2884491.652	;
Input[	316	]=	2728598.85	;
Input[	317	]=	2572463.678	;
Input[	318	]=	2416100.005	;
Input[	319	]=	2259521.72	;
Input[	320	]=	2102742.731	;
Input[	321	]=	1945776.965	;
Input[	322	]=	1788638.363	;
Input[	323	]=	1631340.884	;
Input[	324	]=	1473898.5	;
Input[	325	]=	1316325.196	;
Input[	326	]=	1158634.968	;
Input[	327	]=	1000841.824	;
Input[	328	]=	842959.7789	;
Input[	329	]=	685002.8573	;
Input[	330	]=	526985.0898	;
Input[	331	]=	368920.5124	;
Input[	332	]=	210823.1654	;
Input[	333	]=	52707.09183	;
Input[	334	]=	-105413.6635	;
Input[	335	]=	-263525.0553	;
Input[	336	]=	-421613.0394	;
Input[	337	]=	-579663.5733	;
Input[	338	]=	-737662.6181	;
Input[	339	]=	-895596.1395	;
Input[	340	]=	-1053450.109	;
Input[	341	]=	-1211210.505	;
Input[	342	]=	-1368863.314	;
Input[	343	]=	-1526394.533	;
Input[	344	]=	-1683790.168	;
Input[	345	]=	-1841036.24	;
Input[	346	]=	-1998118.78	;
Input[	347	]=	-2155023.836	;
Input[	348	]=	-2311737.47	;
Input[	349	]=	-2468245.762	;
Input[	350	]=	-2624534.81	;
Input[	351	]=	-2780590.732	;
Input[	352	]=	-2936399.665	;
Input[	353	]=	-3091947.771	;
Input[	354	]=	-3247221.232	;
Input[	355	]=	-3402206.256	;
Input[	356	]=	-3556889.077	;
Input[	357	]=	-3711255.954	;
Input[	358	]=	-3865293.175	;
Input[	359	]=	-4018987.06	;
Input[	360	]=	-4172323.954	;
Input[	361	]=	-4325290.238	;
Input[	362	]=	-4477872.326	;
Input[	363	]=	-4630056.662	;
Input[	364	]=	-4781829.731	;
Input[	365	]=	-4933178.049	;
Input[	366	]=	-5084088.174	;
Input[	367	]=	-5234546.701	;
Input[	368	]=	-5384540.266	;
Input[	369	]=	-5534055.544	;
Input[	370	]=	-5683079.255	;
Input[	371	]=	-5831598.163	;
Input[	372	]=	-5979599.074	;
Input[	373	]=	-6127068.843	;
Input[	374	]=	-6273994.37	;
Input[	375	]=	-6420362.604	;
Input[	376	]=	-6566160.545	;
Input[	377	]=	-6711375.242	;
Input[	378	]=	-6855993.795	;
Input[	379	]=	-7000003.359	;
Input[	380	]=	-7143391.143	;
Input[	381	]=	-7286144.409	;
Input[	382	]=	-7428250.478	;
Input[	383	]=	-7569696.727	;
Input[	384	]=	-7710470.591	;
Input[	385	]=	-7850559.567	;
Input[	386	]=	-7989951.21	;
Input[	387	]=	-8128633.14	;
Input[	388	]=	-8266593.038	;
Input[	389	]=	-8403818.65	;
Input[	390	]=	-8540297.785	;
Input[	391	]=	-8676018.322	;
Input[	392	]=	-8810968.205	;
Input[	393	]=	-8945135.446	;
Input[	394	]=	-9078508.129	;
Input[	395	]=	-9211074.406	;
Input[	396	]=	-9342822.503	;
Input[	397	]=	-9473740.716	;
Input[	398	]=	-9603817.416	;
Input[	399	]=	-9733041.05	;
Input[	400	]=	-9861400.139	;
Input[	401	]=	-9988883.282	;
Input[	402	]=	-10115479.15	;
Input[	403	]=	-10241176.51	;
Input[	404	]=	-10365964.19	;
Input[	405	]=	-10489831.1	;
Input[	406	]=	-10612766.24	;
Input[	407	]=	-10734758.7	;
Input[	408	]=	-10855797.63	;
Input[	409	]=	-10975872.29	;
Input[	410	]=	-11094972.01	;
Input[	411	]=	-11213086.21	;
Input[	412	]=	-11330204.39	;
Input[	413	]=	-11446316.17	;
Input[	414	]=	-11561411.21	;
Input[	415	]=	-11675479.31	;
Input[	416	]=	-11788510.32	;
Input[	417	]=	-11900494.2	;
Input[	418	]=	-12011421.02	;
Input[	419	]=	-12121280.91	;
Input[	420	]=	-12230064.12	;
Input[	421	]=	-12337760.98	;
Input[	422	]=	-12444361.94	;
Input[	423	]=	-12549857.51	;
Input[	424	]=	-12654238.33	;
Input[	425	]=	-12757495.13	;
Input[	426	]=	-12859618.74	;
Input[	427	]=	-12960600.08	;
Input[	428	]=	-13060430.18	;
Input[	429	]=	-13159100.18	;
Input[	430	]=	-13256601.32	;
Input[	431	]=	-13352924.92	;
Input[	432	]=	-13448062.44	;
Input[	433	]=	-13542005.43	;
Input[	434	]=	-13634745.54	;
Input[	435	]=	-13726274.53	;
Input[	436	]=	-13816584.27	;
Input[	437	]=	-13905666.75	;
Input[	438	]=	-13993514.04	;
Input[	439	]=	-14080118.35	;
Input[	440	]=	-14165471.98	;
Input[	441	]=	-14249567.35	;
Input[	442	]=	-14332397	;
Input[	443	]=	-14413953.55	;
Input[	444	]=	-14494229.78	;
Input[	445	]=	-14573218.54	;
Input[	446	]=	-14650912.83	;
Input[	447	]=	-14727305.74	;
Input[	448	]=	-14802390.48	;
Input[	449	]=	-14876160.39	;
Input[	450	]=	-14948608.91	;
Input[	451	]=	-15019729.62	;
Input[	452	]=	-15089516.18	;
Input[	453	]=	-15157962.4	;
Input[	454	]=	-15225062.21	;
Input[	455	]=	-15290809.64	;
Input[	456	]=	-15355198.85	;
Input[	457	]=	-15418224.12	;
Input[	458	]=	-15479879.85	;
Input[	459	]=	-15540160.58	;
Input[	460	]=	-15599060.94	;
Input[	461	]=	-15656575.69	;
Input[	462	]=	-15712699.74	;
Input[	463	]=	-15767428.1	;
Input[	464	]=	-15820755.91	;
Input[	465	]=	-15872678.42	;
Input[	466	]=	-15923191.03	;
Input[	467	]=	-15972289.25	;
Input[	468	]=	-16019968.72	;
Input[	469	]=	-16066225.2	;
Input[	470	]=	-16111054.59	;
Input[	471	]=	-16154452.9	;
Input[	472	]=	-16196416.28	;
Input[	473	]=	-16236941	;
Input[	474	]=	-16276023.46	;
Input[	475	]=	-16313660.19	;
Input[	476	]=	-16349847.84	;
Input[	477	]=	-16384583.21	;
Input[	478	]=	-16417863.21	;
Input[	479	]=	-16449684.87	;
Input[	480	]=	-16480045.38	;
Input[	481	]=	-16508942.04	;
Input[	482	]=	-16536372.27	;
Input[	483	]=	-16562333.65	;
Input[	484	]=	-16586823.87	;
Input[	485	]=	-16609840.75	;
Input[	486	]=	-16631382.25	;
Input[	487	]=	-16651446.45	;
Input[	488	]=	-16670031.58	;
Input[	489	]=	-16687135.97	;
Input[	490	]=	-16702758.12	;
Input[	491	]=	-16716896.63	;
Input[	492	]=	-16729550.26	;
Input[	493	]=	-16740717.86	;
Input[	494	]=	-16750398.46	;
Input[	495	]=	-16758591.19	;
Input[	496	]=	-16765295.33	;
Input[	497	]=	-16770510.28	;
Input[	498	]=	-16774235.57	;
Input[	499	]=	-16776470.88	;
Input[	500	]=	-16777216	;
Input[	501	]=	-16776470.88	;
Input[	502	]=	-16774235.57	;
Input[	503	]=	-16770510.28	;
Input[	504	]=	-16765295.33	;
Input[	505	]=	-16758591.19	;
Input[	506	]=	-16750398.46	;
Input[	507	]=	-16740717.86	;
Input[	508	]=	-16729550.26	;
Input[	509	]=	-16716896.63	;
Input[	510	]=	-16702758.12	;
Input[	511	]=	-16687135.97	;
Input[	512	]=	-16670031.58	;
Input[	513	]=	-16651446.45	;
Input[	514	]=	-16631382.25	;
Input[	515	]=	-16609840.75	;
Input[	516	]=	-16586823.87	;
Input[	517	]=	-16562333.65	;
Input[	518	]=	-16536372.27	;
Input[	519	]=	-16508942.04	;
Input[	520	]=	-16480045.38	;
Input[	521	]=	-16449684.87	;
Input[	522	]=	-16417863.21	;
Input[	523	]=	-16384583.21	;
Input[	524	]=	-16349847.84	;
Input[	525	]=	-16313660.19	;
Input[	526	]=	-16276023.46	;
Input[	527	]=	-16236941	;
Input[	528	]=	-16196416.28	;
Input[	529	]=	-16154452.9	;
Input[	530	]=	-16111054.59	;
Input[	531	]=	-16066225.2	;
Input[	532	]=	-16019968.72	;
Input[	533	]=	-15972289.25	;
Input[	534	]=	-15923191.03	;
Input[	535	]=	-15872678.42	;
Input[	536	]=	-15820755.91	;
Input[	537	]=	-15767428.1	;
Input[	538	]=	-15712699.74	;
Input[	539	]=	-15656575.69	;
Input[	540	]=	-15599060.94	;
Input[	541	]=	-15540160.58	;
Input[	542	]=	-15479879.85	;
Input[	543	]=	-15418224.12	;
Input[	544	]=	-15355198.85	;
Input[	545	]=	-15290809.64	;
Input[	546	]=	-15225062.21	;
Input[	547	]=	-15157962.4	;
Input[	548	]=	-15089516.18	;
Input[	549	]=	-15019729.62	;
Input[	550	]=	-14948608.91	;
Input[	551	]=	-14876160.39	;
Input[	552	]=	-14802390.48	;
Input[	553	]=	-14727305.74	;
Input[	554	]=	-14650912.83	;
Input[	555	]=	-14573218.54	;
Input[	556	]=	-14494229.78	;
Input[	557	]=	-14413953.55	;
Input[	558	]=	-14332397	;
Input[	559	]=	-14249567.35	;
Input[	560	]=	-14165471.98	;
Input[	561	]=	-14080118.35	;
Input[	562	]=	-13993514.04	;
Input[	563	]=	-13905666.75	;
Input[	564	]=	-13816584.27	;
Input[	565	]=	-13726274.53	;
Input[	566	]=	-13634745.54	;
Input[	567	]=	-13542005.43	;
Input[	568	]=	-13448062.44	;
Input[	569	]=	-13352924.92	;
Input[	570	]=	-13256601.32	;
Input[	571	]=	-13159100.18	;
Input[	572	]=	-13060430.18	;
Input[	573	]=	-12960600.08	;
Input[	574	]=	-12859618.74	;
Input[	575	]=	-12757495.13	;
Input[	576	]=	-12654238.33	;
Input[	577	]=	-12549857.51	;
Input[	578	]=	-12444361.94	;
Input[	579	]=	-12337760.98	;
Input[	580	]=	-12230064.12	;
Input[	581	]=	-12121280.91	;
Input[	582	]=	-12011421.02	;
Input[	583	]=	-11900494.2	;
Input[	584	]=	-11788510.32	;
Input[	585	]=	-11675479.31	;
Input[	586	]=	-11561411.21	;
Input[	587	]=	-11446316.17	;
Input[	588	]=	-11330204.39	;
Input[	589	]=	-11213086.21	;
Input[	590	]=	-11094972.01	;
Input[	591	]=	-10975872.29	;
Input[	592	]=	-10855797.63	;
Input[	593	]=	-10734758.7	;
Input[	594	]=	-10612766.24	;
Input[	595	]=	-10489831.1	;
Input[	596	]=	-10365964.19	;
Input[	597	]=	-10241176.51	;
Input[	598	]=	-10115479.15	;
Input[	599	]=	-9988883.282	;
Input[	600	]=	-9861400.139	;
Input[	601	]=	-9733041.05	;
Input[	602	]=	-9603817.416	;
Input[	603	]=	-9473740.716	;
Input[	604	]=	-9342822.503	;
Input[	605	]=	-9211074.406	;
Input[	606	]=	-9078508.129	;
Input[	607	]=	-8945135.446	;
Input[	608	]=	-8810968.205	;
Input[	609	]=	-8676018.322	;
Input[	610	]=	-8540297.785	;
Input[	611	]=	-8403818.65	;
Input[	612	]=	-8266593.038	;
Input[	613	]=	-8128633.14	;
Input[	614	]=	-7989951.21	;
Input[	615	]=	-7850559.567	;
Input[	616	]=	-7710470.591	;
Input[	617	]=	-7569696.727	;
Input[	618	]=	-7428250.478	;
Input[	619	]=	-7286144.409	;
Input[	620	]=	-7143391.143	;
Input[	621	]=	-7000003.359	;
Input[	622	]=	-6855993.795	;
Input[	623	]=	-6711375.242	;
Input[	624	]=	-6566160.545	;
Input[	625	]=	-6420362.604	;
Input[	626	]=	-6273994.37	;
Input[	627	]=	-6127068.843	;
Input[	628	]=	-5979599.074	;
Input[	629	]=	-5831598.163	;
Input[	630	]=	-5683079.255	;
Input[	631	]=	-5534055.544	;
Input[	632	]=	-5384540.266	;
Input[	633	]=	-5234546.701	;
Input[	634	]=	-5084088.174	;
Input[	635	]=	-4933178.049	;
Input[	636	]=	-4781829.731	;
Input[	637	]=	-4630056.662	;
Input[	638	]=	-4477872.326	;
Input[	639	]=	-4325290.238	;
Input[	640	]=	-4172323.954	;
Input[	641	]=	-4018987.06	;
Input[	642	]=	-3865293.175	;
Input[	643	]=	-3711255.954	;
Input[	644	]=	-3556889.077	;
Input[	645	]=	-3402206.256	;
Input[	646	]=	-3247221.232	;
Input[	647	]=	-3091947.771	;
Input[	648	]=	-2936399.665	;
Input[	649	]=	-2780590.732	;
Input[	650	]=	-2624534.81	;
Input[	651	]=	-2468245.762	;
Input[	652	]=	-2311737.47	;
Input[	653	]=	-2155023.836	;
Input[	654	]=	-1998118.78	;
Input[	655	]=	-1841036.24	;
Input[	656	]=	-1683790.168	;
Input[	657	]=	-1526394.533	;
Input[	658	]=	-1368863.314	;
Input[	659	]=	-1211210.505	;
Input[	660	]=	-1053450.109	;
Input[	661	]=	-895596.1395	;
Input[	662	]=	-737662.6181	;
Input[	663	]=	-579663.5733	;
Input[	664	]=	-421613.0394	;
Input[	665	]=	-263525.0553	;
Input[	666	]=	-105413.6635	;

// Tri F = .15 T = .01
//Input[	0	]=	-8388608	;
//Input[	1	]=	-8338276.352	;
//Input[	2	]=	-8287944.704	;
//Input[	3	]=	-8237613.056	;
//Input[	4	]=	-8187281.408	;
//Input[	5	]=	-8136949.76	;
//Input[	6	]=	-8086618.112	;
//Input[	7	]=	-8036286.464	;
//Input[	8	]=	-7985954.816	;
//Input[	9	]=	-7935623.168	;
//Input[	10	]=	-7885291.52	;
//Input[	11	]=	-7834959.872	;
//Input[	12	]=	-7784628.224	;
//Input[	13	]=	-7734296.576	;
//Input[	14	]=	-7683964.928	;
//Input[	15	]=	-7633633.28	;
//Input[	16	]=	-7583301.632	;
//Input[	17	]=	-7532969.984	;
//Input[	18	]=	-7482638.336	;
//Input[	19	]=	-7432306.688	;
//Input[	20	]=	-7381975.04	;
//Input[	21	]=	-7331643.392	;
//Input[	22	]=	-7281311.744	;
//Input[	23	]=	-7230980.096	;
//Input[	24	]=	-7180648.448	;
//Input[	25	]=	-7130316.8	;
//Input[	26	]=	-7079985.152	;
//Input[	27	]=	-7029653.504	;
//Input[	28	]=	-6979321.856	;
//Input[	29	]=	-6928990.208	;
//Input[	30	]=	-6878658.56	;
//Input[	31	]=	-6828326.912	;
//Input[	32	]=	-6777995.264	;
//Input[	33	]=	-6727663.616	;
//Input[	34	]=	-6677331.968	;
//Input[	35	]=	-6627000.32	;
//Input[	36	]=	-6576668.672	;
//Input[	37	]=	-6526337.024	;
//Input[	38	]=	-6476005.376	;
//Input[	39	]=	-6425673.728	;
//Input[	40	]=	-6375342.08	;
//Input[	41	]=	-6325010.432	;
//Input[	42	]=	-6274678.784	;
//Input[	43	]=	-6224347.136	;
//Input[	44	]=	-6174015.488	;
//Input[	45	]=	-6123683.84	;
//Input[	46	]=	-6073352.192	;
//Input[	47	]=	-6023020.544	;
//Input[	48	]=	-5972688.896	;
//Input[	49	]=	-5922357.248	;
//Input[	50	]=	-5872025.6	;
//Input[	51	]=	-5821693.952	;
//Input[	52	]=	-5771362.304	;
//Input[	53	]=	-5721030.656	;
//Input[	54	]=	-5670699.008	;
//Input[	55	]=	-5620367.36	;
//Input[	56	]=	-5570035.712	;
//Input[	57	]=	-5519704.064	;
//Input[	58	]=	-5469372.416	;
//Input[	59	]=	-5419040.768	;
//Input[	60	]=	-5368709.12	;
//Input[	61	]=	-5318377.472	;
//Input[	62	]=	-5268045.824	;
//Input[	63	]=	-5217714.176	;
//Input[	64	]=	-5167382.528	;
//Input[	65	]=	-5117050.88	;
//Input[	66	]=	-5066719.232	;
//Input[	67	]=	-5016387.584	;
//Input[	68	]=	-4966055.936	;
//Input[	69	]=	-4915724.288	;
//Input[	70	]=	-4865392.64	;
//Input[	71	]=	-4815060.992	;
//Input[	72	]=	-4764729.344	;
//Input[	73	]=	-4714397.696	;
//Input[	74	]=	-4664066.048	;
//Input[	75	]=	-4613734.4	;
//Input[	76	]=	-4563402.752	;
//Input[	77	]=	-4513071.104	;
//Input[	78	]=	-4462739.456	;
//Input[	79	]=	-4412407.808	;
//Input[	80	]=	-4362076.16	;
//Input[	81	]=	-4311744.512	;
//Input[	82	]=	-4261412.864	;
//Input[	83	]=	-4211081.216	;
//Input[	84	]=	-4160749.568	;
//Input[	85	]=	-4110417.92	;
//Input[	86	]=	-4060086.272	;
//Input[	87	]=	-4009754.624	;
//Input[	88	]=	-3959422.976	;
//Input[	89	]=	-3909091.328	;
//Input[	90	]=	-3858759.68	;
//Input[	91	]=	-3808428.032	;
//Input[	92	]=	-3758096.384	;
//Input[	93	]=	-3707764.736	;
//Input[	94	]=	-3657433.088	;
//Input[	95	]=	-3607101.44	;
//Input[	96	]=	-3556769.792	;
//Input[	97	]=	-3506438.144	;
//Input[	98	]=	-3456106.496	;
//Input[	99	]=	-3405774.848	;
//Input[	100	]=	-3355443.2	;
//Input[	101	]=	-3305111.552	;
//Input[	102	]=	-3254779.904	;
//Input[	103	]=	-3204448.256	;
//Input[	104	]=	-3154116.608	;
//Input[	105	]=	-3103784.96	;
//Input[	106	]=	-3053453.312	;
//Input[	107	]=	-3003121.664	;
//Input[	108	]=	-2952790.016	;
//Input[	109	]=	-2902458.368	;
//Input[	110	]=	-2852126.72	;
//Input[	111	]=	-2801795.072	;
//Input[	112	]=	-2751463.424	;
//Input[	113	]=	-2701131.776	;
//Input[	114	]=	-2650800.128	;
//Input[	115	]=	-2600468.48	;
//Input[	116	]=	-2550136.832	;
//Input[	117	]=	-2499805.184	;
//Input[	118	]=	-2449473.536	;
//Input[	119	]=	-2399141.888	;
//Input[	120	]=	-2348810.24	;
//Input[	121	]=	-2298478.592	;
//Input[	122	]=	-2248146.944	;
//Input[	123	]=	-2197815.296	;
//Input[	124	]=	-2147483.648	;
//Input[	125	]=	-2097152	;
//Input[	126	]=	-2046820.352	;
//Input[	127	]=	-1996488.704	;
//Input[	128	]=	-1946157.056	;
//Input[	129	]=	-1895825.408	;
//Input[	130	]=	-1845493.76	;
//Input[	131	]=	-1795162.112	;
//Input[	132	]=	-1744830.464	;
//Input[	133	]=	-1694498.816	;
//Input[	134	]=	-1644167.168	;
//Input[	135	]=	-1593835.52	;
//Input[	136	]=	-1543503.872	;
//Input[	137	]=	-1493172.224	;
//Input[	138	]=	-1442840.576	;
//Input[	139	]=	-1392508.928	;
//Input[	140	]=	-1342177.28	;
//Input[	141	]=	-1291845.632	;
//Input[	142	]=	-1241513.984	;
//Input[	143	]=	-1191182.336	;
//Input[	144	]=	-1140850.688	;
//Input[	145	]=	-1090519.04	;
//Input[	146	]=	-1040187.392	;
//Input[	147	]=	-989855.744	;
//Input[	148	]=	-939524.096	;
//Input[	149	]=	-889192.448	;
//Input[	150	]=	-838860.8	;
//Input[	151	]=	-788529.152	;
//Input[	152	]=	-738197.504	;
//Input[	153	]=	-687865.856	;
//Input[	154	]=	-637534.208	;
//Input[	155	]=	-587202.56	;
//Input[	156	]=	-536870.912	;
//Input[	157	]=	-486539.264	;
//Input[	158	]=	-436207.616	;
//Input[	159	]=	-385875.968	;
//Input[	160	]=	-335544.32	;
//Input[	161	]=	-285212.672	;
//Input[	162	]=	-234881.024	;
//Input[	163	]=	-184549.376	;
//Input[	164	]=	-134217.728	;
//Input[	165	]=	-83886.08	;
//Input[	166	]=	-33554.432	;
//Input[	167	]=	16777.216	;
//Input[	168	]=	67108.864	;
//Input[	169	]=	117440.512	;
//Input[	170	]=	167772.16	;
//Input[	171	]=	218103.808	;
//Input[	172	]=	268435.456	;
//Input[	173	]=	318767.104	;
//Input[	174	]=	369098.752	;
//Input[	175	]=	419430.4	;
//Input[	176	]=	469762.048	;
//Input[	177	]=	520093.696	;
//Input[	178	]=	570425.344	;
//Input[	179	]=	620756.992	;
//Input[	180	]=	671088.64	;
//Input[	181	]=	721420.288	;
//Input[	182	]=	771751.936	;
//Input[	183	]=	822083.584	;
//Input[	184	]=	872415.232	;
//Input[	185	]=	922746.88	;
//Input[	186	]=	973078.528	;
//Input[	187	]=	1023410.176	;
//Input[	188	]=	1073741.824	;
//Input[	189	]=	1124073.472	;
//Input[	190	]=	1174405.12	;
//Input[	191	]=	1224736.768	;
//Input[	192	]=	1275068.416	;
//Input[	193	]=	1325400.064	;
//Input[	194	]=	1375731.712	;
//Input[	195	]=	1426063.36	;
//Input[	196	]=	1476395.008	;
//Input[	197	]=	1526726.656	;
//Input[	198	]=	1577058.304	;
//Input[	199	]=	1627389.952	;
//Input[	200	]=	1677721.6	;
//Input[	201	]=	1728053.248	;
//Input[	202	]=	1778384.896	;
//Input[	203	]=	1828716.544	;
//Input[	204	]=	1879048.192	;
//Input[	205	]=	1929379.84	;
//Input[	206	]=	1979711.488	;
//Input[	207	]=	2030043.136	;
//Input[	208	]=	2080374.784	;
//Input[	209	]=	2130706.432	;
//Input[	210	]=	2181038.08	;
//Input[	211	]=	2231369.728	;
//Input[	212	]=	2281701.376	;
//Input[	213	]=	2332033.024	;
//Input[	214	]=	2382364.672	;
//Input[	215	]=	2432696.32	;
//Input[	216	]=	2483027.968	;
//Input[	217	]=	2533359.616	;
//Input[	218	]=	2583691.264	;
//Input[	219	]=	2634022.912	;
//Input[	220	]=	2684354.56	;
//Input[	221	]=	2734686.208	;
//Input[	222	]=	2785017.856	;
//Input[	223	]=	2835349.504	;
//Input[	224	]=	2885681.152	;
//Input[	225	]=	2936012.8	;
//Input[	226	]=	2986344.448	;
//Input[	227	]=	3036676.096	;
//Input[	228	]=	3087007.744	;
//Input[	229	]=	3137339.392	;
//Input[	230	]=	3187671.04	;
//Input[	231	]=	3238002.688	;
//Input[	232	]=	3288334.336	;
//Input[	233	]=	3338665.984	;
//Input[	234	]=	3388997.632	;
//Input[	235	]=	3439329.28	;
//Input[	236	]=	3489660.928	;
//Input[	237	]=	3539992.576	;
//Input[	238	]=	3590324.224	;
//Input[	239	]=	3640655.872	;
//Input[	240	]=	3690987.52	;
//Input[	241	]=	3741319.168	;
//Input[	242	]=	3791650.816	;
//Input[	243	]=	3841982.464	;
//Input[	244	]=	3892314.112	;
//Input[	245	]=	3942645.76	;
//Input[	246	]=	3992977.408	;
//Input[	247	]=	4043309.056	;
//Input[	248	]=	4093640.704	;
//Input[	249	]=	4143972.352	;
//Input[	250	]=	4194304	;
//Input[	251	]=	4244635.648	;
//Input[	252	]=	4294967.296	;
//Input[	253	]=	4345298.944	;
//Input[	254	]=	4395630.592	;
//Input[	255	]=	4445962.24	;
//Input[	256	]=	4496293.888	;
//Input[	257	]=	4546625.536	;
//Input[	258	]=	4596957.184	;
//Input[	259	]=	4647288.832	;
//Input[	260	]=	4697620.48	;
//Input[	261	]=	4747952.128	;
//Input[	262	]=	4798283.776	;
//Input[	263	]=	4848615.424	;
//Input[	264	]=	4898947.072	;
//Input[	265	]=	4949278.72	;
//Input[	266	]=	4999610.368	;
//Input[	267	]=	5049942.016	;
//Input[	268	]=	5100273.664	;
//Input[	269	]=	5150605.312	;
//Input[	270	]=	5200936.96	;
//Input[	271	]=	5251268.608	;
//Input[	272	]=	5301600.256	;
//Input[	273	]=	5351931.904	;
//Input[	274	]=	5402263.552	;
//Input[	275	]=	5452595.2	;
//Input[	276	]=	5502926.848	;
//Input[	277	]=	5553258.496	;
//Input[	278	]=	5603590.144	;
//Input[	279	]=	5653921.792	;
//Input[	280	]=	5704253.44	;
//Input[	281	]=	5754585.088	;
//Input[	282	]=	5804916.736	;
//Input[	283	]=	5855248.384	;
//Input[	284	]=	5905580.032	;
//Input[	285	]=	5955911.68	;
//Input[	286	]=	6006243.328	;
//Input[	287	]=	6056574.976	;
//Input[	288	]=	6106906.624	;
//Input[	289	]=	6157238.272	;
//Input[	290	]=	6207569.92	;
//Input[	291	]=	6257901.568	;
//Input[	292	]=	6308233.216	;
//Input[	293	]=	6358564.864	;
//Input[	294	]=	6408896.512	;
//Input[	295	]=	6459228.16	;
//Input[	296	]=	6509559.808	;
//Input[	297	]=	6559891.456	;
//Input[	298	]=	6610223.104	;
//Input[	299	]=	6660554.752	;
//Input[	300	]=	6710886.4	;
//Input[	301	]=	6761218.048	;
//Input[	302	]=	6811549.696	;
//Input[	303	]=	6861881.344	;
//Input[	304	]=	6912212.992	;
//Input[	305	]=	6962544.64	;
//Input[	306	]=	7012876.288	;
//Input[	307	]=	7063207.936	;
//Input[	308	]=	7113539.584	;
//Input[	309	]=	7163871.232	;
//Input[	310	]=	7214202.88	;
//Input[	311	]=	7264534.528	;
//Input[	312	]=	7314866.176	;
//Input[	313	]=	7365197.824	;
//Input[	314	]=	7415529.472	;
//Input[	315	]=	7465861.12	;
//Input[	316	]=	7516192.768	;
//Input[	317	]=	7566524.416	;
//Input[	318	]=	7616856.064	;
//Input[	319	]=	7667187.712	;
//Input[	320	]=	7717519.36	;
//Input[	321	]=	7767851.008	;
//Input[	322	]=	7818182.656	;
//Input[	323	]=	7868514.304	;
//Input[	324	]=	7918845.952	;
//Input[	325	]=	7969177.6	;
//Input[	326	]=	8019509.248	;
//Input[	327	]=	8069840.896	;
//Input[	328	]=	8120172.544	;
//Input[	329	]=	8170504.192	;
//Input[	330	]=	8220835.84	;
//Input[	331	]=	8271167.488	;
//Input[	332	]=	8321499.136	;
//Input[	333	]=	8371830.784	;
//Input[	334	]=	8355053.568	;
//Input[	335	]=	8304721.92	;
//Input[	336	]=	8254390.272	;
//Input[	337	]=	8204058.624	;
//Input[	338	]=	8153726.976	;
//Input[	339	]=	8103395.328	;
//Input[	340	]=	8053063.68	;
//Input[	341	]=	8002732.032	;
//Input[	342	]=	7952400.384	;
//Input[	343	]=	7902068.736	;
//Input[	344	]=	7851737.088	;
//Input[	345	]=	7801405.44	;
//Input[	346	]=	7751073.792	;
//Input[	347	]=	7700742.144	;
//Input[	348	]=	7650410.496	;
//Input[	349	]=	7600078.848	;
//Input[	350	]=	7549747.2	;
//Input[	351	]=	7499415.552	;
//Input[	352	]=	7449083.904	;
//Input[	353	]=	7398752.256	;
//Input[	354	]=	7348420.608	;
//Input[	355	]=	7298088.96	;
//Input[	356	]=	7247757.312	;
//Input[	357	]=	7197425.664	;
//Input[	358	]=	7147094.016	;
//Input[	359	]=	7096762.368	;
//Input[	360	]=	7046430.72	;
//Input[	361	]=	6996099.072	;
//Input[	362	]=	6945767.424	;
//Input[	363	]=	6895435.776	;
//Input[	364	]=	6845104.128	;
//Input[	365	]=	6794772.48	;
//Input[	366	]=	6744440.832	;
//Input[	367	]=	6694109.184	;
//Input[	368	]=	6643777.536	;
//Input[	369	]=	6593445.888	;
//Input[	370	]=	6543114.24	;
//Input[	371	]=	6492782.592	;
//Input[	372	]=	6442450.944	;
//Input[	373	]=	6392119.296	;
//Input[	374	]=	6341787.648	;
//Input[	375	]=	6291456	;
//Input[	376	]=	6241124.352	;
//Input[	377	]=	6190792.704	;
//Input[	378	]=	6140461.056	;
//Input[	379	]=	6090129.408	;
//Input[	380	]=	6039797.76	;
//Input[	381	]=	5989466.112	;
//Input[	382	]=	5939134.464	;
//Input[	383	]=	5888802.816	;
//Input[	384	]=	5838471.168	;
//Input[	385	]=	5788139.52	;
//Input[	386	]=	5737807.872	;
//Input[	387	]=	5687476.224	;
//Input[	388	]=	5637144.576	;
//Input[	389	]=	5586812.928	;
//Input[	390	]=	5536481.28	;
//Input[	391	]=	5486149.632	;
//Input[	392	]=	5435817.984	;
//Input[	393	]=	5385486.336	;
//Input[	394	]=	5335154.688	;
//Input[	395	]=	5284823.04	;
//Input[	396	]=	5234491.392	;
//Input[	397	]=	5184159.744	;
//Input[	398	]=	5133828.096	;
//Input[	399	]=	5083496.448	;
//Input[	400	]=	5033164.8	;
//Input[	401	]=	4982833.152	;
//Input[	402	]=	4932501.504	;
//Input[	403	]=	4882169.856	;
//Input[	404	]=	4831838.208	;
//Input[	405	]=	4781506.56	;
//Input[	406	]=	4731174.912	;
//Input[	407	]=	4680843.264	;
//Input[	408	]=	4630511.616	;
//Input[	409	]=	4580179.968	;
//Input[	410	]=	4529848.32	;
//Input[	411	]=	4479516.672	;
//Input[	412	]=	4429185.024	;
//Input[	413	]=	4378853.376	;
//Input[	414	]=	4328521.728	;
//Input[	415	]=	4278190.08	;
//Input[	416	]=	4227858.432	;
//Input[	417	]=	4177526.784	;
//Input[	418	]=	4127195.136	;
//Input[	419	]=	4076863.488	;
//Input[	420	]=	4026531.84	;
//Input[	421	]=	3976200.192	;
//Input[	422	]=	3925868.544	;
//Input[	423	]=	3875536.896	;
//Input[	424	]=	3825205.248	;
//Input[	425	]=	3774873.6	;
//Input[	426	]=	3724541.952	;
//Input[	427	]=	3674210.304	;
//Input[	428	]=	3623878.656	;
//Input[	429	]=	3573547.008	;
//Input[	430	]=	3523215.36	;
//Input[	431	]=	3472883.712	;
//Input[	432	]=	3422552.064	;
//Input[	433	]=	3372220.416	;
//Input[	434	]=	3321888.768	;
//Input[	435	]=	3271557.12	;
//Input[	436	]=	3221225.472	;
//Input[	437	]=	3170893.824	;
//Input[	438	]=	3120562.176	;
//Input[	439	]=	3070230.528	;
//Input[	440	]=	3019898.88	;
//Input[	441	]=	2969567.232	;
//Input[	442	]=	2919235.584	;
//Input[	443	]=	2868903.936	;
//Input[	444	]=	2818572.288	;
//Input[	445	]=	2768240.64	;
//Input[	446	]=	2717908.992	;
//Input[	447	]=	2667577.344	;
//Input[	448	]=	2617245.696	;
//Input[	449	]=	2566914.048	;
//Input[	450	]=	2516582.4	;
//Input[	451	]=	2466250.752	;
//Input[	452	]=	2415919.104	;
//Input[	453	]=	2365587.456	;
//Input[	454	]=	2315255.808	;
//Input[	455	]=	2264924.16	;
//Input[	456	]=	2214592.512	;
//Input[	457	]=	2164260.864	;
//Input[	458	]=	2113929.216	;
//Input[	459	]=	2063597.568	;
//Input[	460	]=	2013265.92	;
//Input[	461	]=	1962934.272	;
//Input[	462	]=	1912602.624	;
//Input[	463	]=	1862270.976	;
//Input[	464	]=	1811939.328	;
//Input[	465	]=	1761607.68	;
//Input[	466	]=	1711276.032	;
//Input[	467	]=	1660944.384	;
//Input[	468	]=	1610612.736	;
//Input[	469	]=	1560281.088	;
//Input[	470	]=	1509949.44	;
//Input[	471	]=	1459617.792	;
//Input[	472	]=	1409286.144	;
//Input[	473	]=	1358954.496	;
//Input[	474	]=	1308622.848	;
//Input[	475	]=	1258291.2	;
//Input[	476	]=	1207959.552	;
//Input[	477	]=	1157627.904	;
//Input[	478	]=	1107296.256	;
//Input[	479	]=	1056964.608	;
//Input[	480	]=	1006632.96	;
//Input[	481	]=	956301.312	;
//Input[	482	]=	905969.664	;
//Input[	483	]=	855638.016	;
//Input[	484	]=	805306.368	;
//Input[	485	]=	754974.72	;
//Input[	486	]=	704643.072	;
//Input[	487	]=	654311.424	;
//Input[	488	]=	603979.776	;
//Input[	489	]=	553648.128	;
//Input[	490	]=	503316.48	;
//Input[	491	]=	452984.832	;
//Input[	492	]=	402653.184	;
//Input[	493	]=	352321.536	;
//Input[	494	]=	301989.888	;
//Input[	495	]=	251658.24	;
//Input[	496	]=	201326.592	;
//Input[	497	]=	150994.944	;
//Input[	498	]=	100663.296	;
//Input[	499	]=	50331.648	;
//Input[	500	]=	0	;
//Input[	501	]=	-50331.648	;
//Input[	502	]=	-100663.296	;
//Input[	503	]=	-150994.944	;
//Input[	504	]=	-201326.592	;
//Input[	505	]=	-251658.24	;
//Input[	506	]=	-301989.888	;
//Input[	507	]=	-352321.536	;
//Input[	508	]=	-402653.184	;
//Input[	509	]=	-452984.832	;
//Input[	510	]=	-503316.48	;
//Input[	511	]=	-553648.128	;
//Input[	512	]=	-603979.776	;
//Input[	513	]=	-654311.424	;
//Input[	514	]=	-704643.072	;
//Input[	515	]=	-754974.72	;
//Input[	516	]=	-805306.368	;
//Input[	517	]=	-855638.016	;
//Input[	518	]=	-905969.664	;
//Input[	519	]=	-956301.312	;
//Input[	520	]=	-1006632.96	;
//Input[	521	]=	-1056964.608	;
//Input[	522	]=	-1107296.256	;
//Input[	523	]=	-1157627.904	;
//Input[	524	]=	-1207959.552	;
//Input[	525	]=	-1258291.2	;
//Input[	526	]=	-1308622.848	;
//Input[	527	]=	-1358954.496	;
//Input[	528	]=	-1409286.144	;
//Input[	529	]=	-1459617.792	;
//Input[	530	]=	-1509949.44	;
//Input[	531	]=	-1560281.088	;
//Input[	532	]=	-1610612.736	;
//Input[	533	]=	-1660944.384	;
//Input[	534	]=	-1711276.032	;
//Input[	535	]=	-1761607.68	;
//Input[	536	]=	-1811939.328	;
//Input[	537	]=	-1862270.976	;
//Input[	538	]=	-1912602.624	;
//Input[	539	]=	-1962934.272	;
//Input[	540	]=	-2013265.92	;
//Input[	541	]=	-2063597.568	;
//Input[	542	]=	-2113929.216	;
//Input[	543	]=	-2164260.864	;
//Input[	544	]=	-2214592.512	;
//Input[	545	]=	-2264924.16	;
//Input[	546	]=	-2315255.808	;
//Input[	547	]=	-2365587.456	;
//Input[	548	]=	-2415919.104	;
//Input[	549	]=	-2466250.752	;
//Input[	550	]=	-2516582.4	;
//Input[	551	]=	-2566914.048	;
//Input[	552	]=	-2617245.696	;
//Input[	553	]=	-2667577.344	;
//Input[	554	]=	-2717908.992	;
//Input[	555	]=	-2768240.64	;
//Input[	556	]=	-2818572.288	;
//Input[	557	]=	-2868903.936	;
//Input[	558	]=	-2919235.584	;
//Input[	559	]=	-2969567.232	;
//Input[	560	]=	-3019898.88	;
//Input[	561	]=	-3070230.528	;
//Input[	562	]=	-3120562.176	;
//Input[	563	]=	-3170893.824	;
//Input[	564	]=	-3221225.472	;
//Input[	565	]=	-3271557.12	;
//Input[	566	]=	-3321888.768	;
//Input[	567	]=	-3372220.416	;
//Input[	568	]=	-3422552.064	;
//Input[	569	]=	-3472883.712	;
//Input[	570	]=	-3523215.36	;
//Input[	571	]=	-3573547.008	;
//Input[	572	]=	-3623878.656	;
//Input[	573	]=	-3674210.304	;
//Input[	574	]=	-3724541.952	;
//Input[	575	]=	-3774873.6	;
//Input[	576	]=	-3825205.248	;
//Input[	577	]=	-3875536.896	;
//Input[	578	]=	-3925868.544	;
//Input[	579	]=	-3976200.192	;
//Input[	580	]=	-4026531.84	;
//Input[	581	]=	-4076863.488	;
//Input[	582	]=	-4127195.136	;
//Input[	583	]=	-4177526.784	;
//Input[	584	]=	-4227858.432	;
//Input[	585	]=	-4278190.08	;
//Input[	586	]=	-4328521.728	;
//Input[	587	]=	-4378853.376	;
//Input[	588	]=	-4429185.024	;
//Input[	589	]=	-4479516.672	;
//Input[	590	]=	-4529848.32	;
//Input[	591	]=	-4580179.968	;
//Input[	592	]=	-4630511.616	;
//Input[	593	]=	-4680843.264	;
//Input[	594	]=	-4731174.912	;
//Input[	595	]=	-4781506.56	;
//Input[	596	]=	-4831838.208	;
//Input[	597	]=	-4882169.856	;
//Input[	598	]=	-4932501.504	;
//Input[	599	]=	-4982833.152	;
//Input[	600	]=	-5033164.8	;
//Input[	601	]=	-5083496.448	;
//Input[	602	]=	-5133828.096	;
//Input[	603	]=	-5184159.744	;
//Input[	604	]=	-5234491.392	;
//Input[	605	]=	-5284823.04	;
//Input[	606	]=	-5335154.688	;
//Input[	607	]=	-5385486.336	;
//Input[	608	]=	-5435817.984	;
//Input[	609	]=	-5486149.632	;
//Input[	610	]=	-5536481.28	;
//Input[	611	]=	-5586812.928	;
//Input[	612	]=	-5637144.576	;
//Input[	613	]=	-5687476.224	;
//Input[	614	]=	-5737807.872	;
//Input[	615	]=	-5788139.52	;
//Input[	616	]=	-5838471.168	;
//Input[	617	]=	-5888802.816	;
//Input[	618	]=	-5939134.464	;
//Input[	619	]=	-5989466.112	;
//Input[	620	]=	-6039797.76	;
//Input[	621	]=	-6090129.408	;
//Input[	622	]=	-6140461.056	;
//Input[	623	]=	-6190792.704	;
//Input[	624	]=	-6241124.352	;
//Input[	625	]=	-6291456	;
//Input[	626	]=	-6341787.648	;
//Input[	627	]=	-6392119.296	;
//Input[	628	]=	-6442450.944	;
//Input[	629	]=	-6492782.592	;
//Input[	630	]=	-6543114.24	;
//Input[	631	]=	-6593445.888	;
//Input[	632	]=	-6643777.536	;
//Input[	633	]=	-6694109.184	;
//Input[	634	]=	-6744440.832	;
//Input[	635	]=	-6794772.48	;
//Input[	636	]=	-6845104.128	;
//Input[	637	]=	-6895435.776	;
//Input[	638	]=	-6945767.424	;
//Input[	639	]=	-6996099.072	;
//Input[	640	]=	-7046430.72	;
//Input[	641	]=	-7096762.368	;
//Input[	642	]=	-7147094.016	;
//Input[	643	]=	-7197425.664	;
//Input[	644	]=	-7247757.312	;
//Input[	645	]=	-7298088.96	;
//Input[	646	]=	-7348420.608	;
//Input[	647	]=	-7398752.256	;
//Input[	648	]=	-7449083.904	;
//Input[	649	]=	-7499415.552	;
//Input[	650	]=	-7549747.2	;
//Input[	651	]=	-7600078.848	;
//Input[	652	]=	-7650410.496	;
//Input[	653	]=	-7700742.144	;
//Input[	654	]=	-7751073.792	;
//Input[	655	]=	-7801405.44	;
//Input[	656	]=	-7851737.088	;
//Input[	657	]=	-7902068.736	;
//Input[	658	]=	-7952400.384	;
//Input[	659	]=	-8002732.032	;
//Input[	660	]=	-8053063.68	;
//Input[	661	]=	-8103395.328	;
//Input[	662	]=	-8153726.976	;
//Input[	663	]=	-8204058.624	;
//Input[	664	]=	-8254390.272	;
//Input[	665	]=	-8304721.92	;
//Input[	666	]=	-8355053.568	;

Signal<=0;
SigInd <=0;

end

always @( posedge control )
begin
	// Output = stored values
	
	
		Signal = Input[i];
		i=i+1;
		SigInd = !SigInd;
		if (i>SigLength)
		begin
		i=0;
		end
end

endmodule
