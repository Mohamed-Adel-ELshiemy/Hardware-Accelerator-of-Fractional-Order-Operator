`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    14:27:11 08/22/2021 
// Design Name: 
// Module Name:    SignalLUT 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module SignalLUT(

	input control,
   input  rst,
	output reg [31:0] Signal,
	output reg SigInd
    );
	
	 
	parameter SignalLength = 1884;
	
	reg signed [31:0] Input [0:SignalLength];
	integer i=0;
initial begin

//////////////////////////////////////////////////////////////////////////////////////////////////////////////////
//////////////////////////////////////////////////////////////////////////////////////////////////////////////////
//// Sawtooth
//Input[0]=-16777216;
//Input[1]=-16723812.4628456;
//Input[2]=-16670408.9256912;
//Input[3]=-16617005.3885368;
//Input[4]=-16563601.8513824;
//Input[5]=-16510198.314228;
//Input[6]=-16456794.7770735;
//Input[7]=-16403391.2399191;
//Input[8]=-16349987.7027647;
//Input[9]=-16296584.1656103;
//Input[10]=-16243180.6284559;
//Input[11]=-16189777.0913015;
//Input[12]=-16136373.5541471;
//Input[13]=-16082970.0169927;
//Input[14]=-16029566.4798383;
//Input[15]=-15976162.9426839;
//Input[16]=-15922759.4055295;
//Input[17]=-15869355.8683751;
//Input[18]=-15815952.3312206;
//Input[19]=-15762548.7940662;
//Input[20]=-15709145.2569118;
//Input[21]=-15655741.7197574;
//Input[22]=-15602338.182603;
//Input[23]=-15548934.6454486;
//Input[24]=-15495531.1082942;
//Input[25]=-15442127.5711398;
//Input[26]=-15388724.0339854;
//Input[27]=-15335320.496831;
//Input[28]=-15281916.9596766;
//Input[29]=-15228513.4225221;
//Input[30]=-15175109.8853677;
//Input[31]=-15121706.3482133;
//Input[32]=-15068302.8110589;
//Input[33]=-15014899.2739045;
//Input[34]=-14961495.7367501;
//Input[35]=-14908092.1995957;
//Input[36]=-14854688.6624413;
//Input[37]=-14801285.1252869;
//Input[38]=-14747881.5881325;
//Input[39]=-14694478.0509781;
//Input[40]=-14641074.5138237;
//Input[41]=-14587670.9766692;
//Input[42]=-14534267.4395148;
//Input[43]=-14480863.9023604;
//Input[44]=-14427460.365206;
//Input[45]=-14374056.8280516;
//Input[46]=-14320653.2908972;
//Input[47]=-14267249.7537428;
//Input[48]=-14213846.2165884;
//Input[49]=-14160442.679434;
//Input[50]=-14107039.1422796;
//Input[51]=-14053635.6051252;
//Input[52]=-14000232.0679707;
//Input[53]=-13946828.5308163;
//Input[54]=-13893424.9936619;
//Input[55]=-13840021.4565075;
//Input[56]=-13786617.9193531;
//Input[57]=-13733214.3821987;
//Input[58]=-13679810.8450443;
//Input[59]=-13626407.3078899;
//Input[60]=-13573003.7707355;
//Input[61]=-13519600.2335811;
//Input[62]=-13466196.6964267;
//Input[63]=-13412793.1592723;
//Input[64]=-13359389.6221178;
//Input[65]=-13305986.0849634;
//Input[66]=-13252582.547809;
//Input[67]=-13199179.0106546;
//Input[68]=-13145775.4735002;
//Input[69]=-13092371.9363458;
//Input[70]=-13038968.3991914;
//Input[71]=-12985564.862037;
//Input[72]=-12932161.3248826;
//Input[73]=-12878757.7877282;
//Input[74]=-12825354.2505738;
//Input[75]=-12771950.7134193;
//Input[76]=-12718547.1762649;
//Input[77]=-12665143.6391105;
//Input[78]=-12611740.1019561;
//Input[79]=-12558336.5648017;
//Input[80]=-12504933.0276473;
//Input[81]=-12451529.4904929;
//Input[82]=-12398125.9533385;
//Input[83]=-12344722.4161841;
//Input[84]=-12291318.8790297;
//Input[85]=-12237915.3418753;
//Input[86]=-12184511.8047208;
//Input[87]=-12131108.2675664;
//Input[88]=-12077704.730412;
//Input[89]=-12024301.1932576;
//Input[90]=-11970897.6561032;
//Input[91]=-11917494.1189488;
//Input[92]=-11864090.5817944;
//Input[93]=-11810687.04464;
//Input[94]=-11757283.5074856;
//Input[95]=-11703879.9703312;
//Input[96]=-11650476.4331768;
//Input[97]=-11597072.8960224;
//Input[98]=-11543669.3588679;
//Input[99]=-11490265.8217135;
//Input[100]=-11436862.2845591;
//Input[101]=-11383458.7474047;
//Input[102]=-11330055.2102503;
//Input[103]=-11276651.6730959;
//Input[104]=-11223248.1359415;
//Input[105]=-11169844.5987871;
//Input[106]=-11116441.0616327;
//Input[107]=-11063037.5244783;
//Input[108]=-11009633.9873239;
//Input[109]=-10956230.4501694;
//Input[110]=-10902826.913015;
//Input[111]=-10849423.3758606;
//Input[112]=-10796019.8387062;
//Input[113]=-10742616.3015518;
//Input[114]=-10689212.7643974;
//Input[115]=-10635809.227243;
//Input[116]=-10582405.6900886;
//Input[117]=-10529002.1529342;
//Input[118]=-10475598.6157798;
//Input[119]=-10422195.0786254;
//Input[120]=-10368791.541471;
//Input[121]=-10315388.0043165;
//Input[122]=-10261984.4671621;
//Input[123]=-10208580.9300077;
//Input[124]=-10155177.3928533;
//Input[125]=-10101773.8556989;
//Input[126]=-10048370.3185445;
//Input[127]=-9994966.78139009;
//Input[128]=-9941563.24423568;
//Input[129]=-9888159.70708128;
//Input[130]=-9834756.16992687;
//Input[131]=-9781352.63277246;
//Input[132]=-9727949.09561805;
//Input[133]=-9674545.55846364;
//Input[134]=-9621142.02130923;
//Input[135]=-9567738.48415482;
//Input[136]=-9514334.94700041;
//Input[137]=-9460931.409846;
//Input[138]=-9407527.8726916;
//Input[139]=-9354124.33553719;
//Input[140]=-9300720.79838278;
//Input[141]=-9247317.26122837;
//Input[142]=-9193913.72407396;
//Input[143]=-9140510.18691955;
//Input[144]=-9087106.64976515;
//Input[145]=-9033703.11261074;
//Input[146]=-8980299.57545633;
//Input[147]=-8926896.03830192;
//Input[148]=-8873492.50114751;
//Input[149]=-8820088.9639931;
//Input[150]=-8766685.42683869;
//Input[151]=-8713281.88968428;
//Input[152]=-8659878.35252987;
//Input[153]=-8606474.81537547;
//Input[154]=-8553071.27822106;
//Input[155]=-8499667.74106665;
//Input[156]=-8446264.20391224;
//Input[157]=-8392860.66675783;
//Input[158]=-8339457.12960342;
//Input[159]=-8286053.59244901;
//Input[160]=-8232650.05529461;
//Input[161]=-8179246.5181402;
//Input[162]=-8125842.98098579;
//Input[163]=-8072439.44383138;
//Input[164]=-8019035.90667697;
//Input[165]=-7965632.36952256;
//Input[166]=-7912228.83236815;
//Input[167]=-7858825.29521374;
//Input[168]=-7805421.75805934;
//Input[169]=-7752018.22090493;
//Input[170]=-7698614.68375052;
//Input[171]=-7645211.14659611;
//Input[172]=-7591807.6094417;
//Input[173]=-7538404.07228729;
//Input[174]=-7485000.53513288;
//Input[175]=-7431596.99797847;
//Input[176]=-7378193.46082407;
//Input[177]=-7324789.92366966;
//Input[178]=-7271386.38651525;
//Input[179]=-7217982.84936084;
//Input[180]=-7164579.31220643;
//Input[181]=-7111175.77505202;
//Input[182]=-7057772.23789761;
//Input[183]=-7004368.7007432;
//Input[184]=-6950965.16358879;
//Input[185]=-6897561.62643439;
//Input[186]=-6844158.08927998;
//Input[187]=-6790754.55212557;
//Input[188]=-6737351.01497116;
//Input[189]=-6683947.47781675;
//Input[190]=-6630543.94066234;
//Input[191]=-6577140.40350793;
//Input[192]=-6523736.86635353;
//Input[193]=-6470333.32919912;
//Input[194]=-6416929.79204471;
//Input[195]=-6363526.2548903;
//Input[196]=-6310122.71773589;
//Input[197]=-6256719.18058148;
//Input[198]=-6203315.64342707;
//Input[199]=-6149912.10627266;
//Input[200]=-6096508.56911826;
//Input[201]=-6043105.03196385;
//Input[202]=-5989701.49480944;
//Input[203]=-5936297.95765503;
//Input[204]=-5882894.42050062;
//Input[205]=-5829490.88334621;
//Input[206]=-5776087.3461918;
//Input[207]=-5722683.8090374;
//Input[208]=-5669280.27188299;
//Input[209]=-5615876.73472858;
//Input[210]=-5562473.19757417;
//Input[211]=-5509069.66041976;
//Input[212]=-5455666.12326535;
//Input[213]=-5402262.58611094;
//Input[214]=-5348859.04895653;
//Input[215]=-5295455.51180213;
//Input[216]=-5242051.97464772;
//Input[217]=-5188648.43749331;
//Input[218]=-5135244.9003389;
//Input[219]=-5081841.36318449;
//Input[220]=-5028437.82603008;
//Input[221]=-4975034.28887567;
//Input[222]=-4921630.75172126;
//Input[223]=-4868227.21456686;
//Input[224]=-4814823.67741245;
//Input[225]=-4761420.14025804;
//Input[226]=-4708016.60310363;
//Input[227]=-4654613.06594922;
//Input[228]=-4601209.52879481;
//Input[229]=-4547805.9916404;
//Input[230]=-4494402.45448599;
//Input[231]=-4440998.91733159;
//Input[232]=-4387595.38017718;
//Input[233]=-4334191.84302277;
//Input[234]=-4280788.30586836;
//Input[235]=-4227384.76871395;
//Input[236]=-4173981.23155954;
//Input[237]=-4120577.69440513;
//Input[238]=-4067174.15725072;
//Input[239]=-4013770.62009631;
//Input[240]=-3960367.08294191;
//Input[241]=-3906963.5457875;
//Input[242]=-3853560.00863309;
//Input[243]=-3800156.47147868;
//Input[244]=-3746752.93432427;
//Input[245]=-3693349.39716986;
//Input[246]=-3639945.86001546;
//Input[247]=-3586542.32286105;
//Input[248]=-3533138.78570664;
//Input[249]=-3479735.24855223;
//Input[250]=-3426331.71139782;
//Input[251]=-3372928.17424341;
//Input[252]=-3319524.637089;
//Input[253]=-3266121.09993459;
//Input[254]=-3212717.56278018;
//Input[255]=-3159314.02562577;
//Input[256]=-3105910.48847137;
//Input[257]=-3052506.95131696;
//Input[258]=-2999103.41416255;
//Input[259]=-2945699.87700814;
//Input[260]=-2892296.33985373;
//Input[261]=-2838892.80269932;
//Input[262]=-2785489.26554491;
//Input[263]=-2732085.72839051;
//Input[264]=-2678682.1912361;
//Input[265]=-2625278.65408169;
//Input[266]=-2571875.11692728;
//Input[267]=-2518471.57977287;
//Input[268]=-2465068.04261846;
//Input[269]=-2411664.50546405;
//Input[270]=-2358260.96830964;
//Input[271]=-2304857.43115524;
//Input[272]=-2251453.89400083;
//Input[273]=-2198050.35684642;
//Input[274]=-2144646.81969201;
//Input[275]=-2091243.2825376;
//Input[276]=-2037839.74538319;
//Input[277]=-1984436.20822878;
//Input[278]=-1931032.67107437;
//Input[279]=-1877629.13391997;
//Input[280]=-1824225.59676556;
//Input[281]=-1770822.05961115;
//Input[282]=-1717418.52245674;
//Input[283]=-1664014.98530233;
//Input[284]=-1610611.44814792;
//Input[285]=-1557207.91099351;
//Input[286]=-1503804.37383911;
//Input[287]=-1450400.8366847;
//Input[288]=-1396997.29953029;
//Input[289]=-1343593.76237588;
//Input[290]=-1290190.22522147;
//Input[291]=-1236786.68806706;
//Input[292]=-1183383.15091265;
//Input[293]=-1129979.61375824;
//Input[294]=-1076576.07660384;
//Input[295]=-1023172.53944943;
//Input[296]=-969769.002295019;
//Input[297]=-916365.465140609;
//Input[298]=-862961.927986201;
//Input[299]=-809558.390831791;
//Input[300]=-756154.853677385;
//Input[301]=-702751.316522975;
//Input[302]=-649347.779368566;
//Input[303]=-595944.242214156;
//Input[304]=-542540.705059748;
//Input[305]=-489137.167905338;
//Input[306]=-435733.630750932;
//Input[307]=-382330.093596522;
//Input[308]=-328926.556442114;
//Input[309]=-275523.019287705;
//Input[310]=-222119.482133295;
//Input[311]=-168715.944978889;
//Input[312]=-115312.407824479;
//Input[313]=-61908.8706700709;
//Input[314]=-8505.33351566084;
//Input[315]=44898.2036387473;
//Input[316]=98301.7407931574;
//Input[317]=151705.277947564;
//Input[318]=205108.815101974;
//Input[319]=258512.35225638;
//Input[320]=311915.88941079;
//Input[321]=365319.4265652;
//Input[322]=418722.96371961;
//Input[323]=472126.500874016;
//Input[324]=525530.038028427;
//Input[325]=578933.575182833;
//Input[326]=632337.112337243;
//Input[327]=685740.649491653;
//Input[328]=739144.186646063;
//Input[329]=792547.723800469;
//Input[330]=845951.260954879;
//Input[331]=899354.798109286;
//Input[332]=952758.335263696;
//Input[333]=1006161.87241811;
//Input[334]=1059565.40957251;
//Input[335]=1112968.94672692;
//Input[336]=1166372.48388133;
//Input[337]=1219776.02103574;
//Input[338]=1273179.55819015;
//Input[339]=1326583.09534456;
//Input[340]=1379986.63249896;
//Input[341]=1433390.16965337;
//Input[342]=1486793.70680778;
//Input[343]=1540197.24396219;
//Input[344]=1593600.7811166;
//Input[345]=1647004.31827101;
//Input[346]=1700407.85542542;
//Input[347]=1753811.39257983;
//Input[348]=1807214.92973423;
//Input[349]=1860618.46688864;
//Input[350]=1914022.00404305;
//Input[351]=1967425.54119746;
//Input[352]=2020829.07835187;
//Input[353]=2074232.61550628;
//Input[354]=2127636.15266069;
//Input[355]=2181039.6898151;
//Input[356]=2234443.22696951;
//Input[357]=2287846.76412392;
//Input[358]=2341250.30127832;
//Input[359]=2394653.83843273;
//Input[360]=2448057.37558714;
//Input[361]=2501460.91274155;
//Input[362]=2554864.44989596;
//Input[363]=2608267.98705037;
//Input[364]=2661671.52420478;
//Input[365]=2715075.06135918;
//Input[366]=2768478.59851359;
//Input[367]=2821882.135668;
//Input[368]=2875285.67282241;
//Input[369]=2928689.20997682;
//Input[370]=2982092.74713123;
//Input[371]=3035496.28428563;
//Input[372]=3088899.82144005;
//Input[373]=3142303.35859445;
//Input[374]=3195706.89574886;
//Input[375]=3249110.43290327;
//Input[376]=3302513.97005768;
//Input[377]=3355917.50721209;
//Input[378]=3409321.0443665;
//Input[379]=3462724.5815209;
//Input[380]=3516128.11867531;
//Input[381]=3569531.65582972;
//Input[382]=3622935.19298413;
//Input[383]=3676338.73013854;
//Input[384]=3729742.26729295;
//Input[385]=3783145.80444736;
//Input[386]=3836549.34160177;
//Input[387]=3889952.87875618;
//Input[388]=3943356.41591058;
//Input[389]=3996759.95306499;
//Input[390]=4050163.4902194;
//Input[391]=4103567.02737381;
//Input[392]=4156970.56452822;
//Input[393]=4210374.10168263;
//Input[394]=4263777.63883704;
//Input[395]=4317181.17599145;
//Input[396]=4370584.71314585;
//Input[397]=4423988.25030026;
//Input[398]=4477391.78745467;
//Input[399]=4530795.32460908;
//Input[400]=4584198.86176349;
//Input[401]=4637602.3989179;
//Input[402]=4691005.93607231;
//Input[403]=4744409.47322672;
//Input[404]=4797813.01038113;
//Input[405]=4851216.54753553;
//Input[406]=4904620.08468995;
//Input[407]=4958023.62184435;
//Input[408]=5011427.15899876;
//Input[409]=5064830.69615317;
//Input[410]=5118234.23330757;
//Input[411]=5171637.77046199;
//Input[412]=5225041.30761639;
//Input[413]=5278444.8447708;
//Input[414]=5331848.38192521;
//Input[415]=5385251.91907962;
//Input[416]=5438655.45623403;
//Input[417]=5492058.99338844;
//Input[418]=5545462.53054284;
//Input[419]=5598866.06769726;
//Input[420]=5652269.60485166;
//Input[421]=5705673.14200607;
//Input[422]=5759076.67916048;
//Input[423]=5812480.21631489;
//Input[424]=5865883.7534693;
//Input[425]=5919287.29062371;
//Input[426]=5972690.82777812;
//Input[427]=6026094.36493253;
//Input[428]=6079497.90208693;
//Input[429]=6132901.43924134;
//Input[430]=6186304.97639575;
//Input[431]=6239708.51355016;
//Input[432]=6293112.05070457;
//Input[433]=6346515.58785898;
//Input[434]=6399919.12501339;
//Input[435]=6453322.6621678;
//Input[436]=6506726.19932221;
//Input[437]=6560129.73647661;
//Input[438]=6613533.27363102;
//Input[439]=6666936.81078543;
//Input[440]=6720340.34793984;
//Input[441]=6773743.88509425;
//Input[442]=6827147.42224865;
//Input[443]=6880550.95940306;
//Input[444]=6933954.49655747;
//Input[445]=6987358.03371188;
//Input[446]=7040761.57086629;
//Input[447]=7094165.1080207;
//Input[448]=7147568.64517511;
//Input[449]=7200972.18232952;
//Input[450]=7254375.71948392;
//Input[451]=7307779.25663833;
//Input[452]=7361182.79379274;
//Input[453]=7414586.33094715;
//Input[454]=7467989.86810156;
//Input[455]=7521393.40525597;
//Input[456]=7574796.94241038;
//Input[457]=7628200.47956479;
//Input[458]=7681604.0167192;
//Input[459]=7735007.5538736;
//Input[460]=7788411.09102802;
//Input[461]=7841814.62818242;
//Input[462]=7895218.16533683;
//Input[463]=7948621.70249124;
//Input[464]=8002025.23964565;
//Input[465]=8055428.77680006;
//Input[466]=8108832.31395447;
//Input[467]=8162235.85110887;
//Input[468]=8215639.38826328;
//Input[469]=8269042.92541769;
//Input[470]=8322446.4625721;
//Input[471]=8375849.99972651;
//Input[472]=8429253.53688091;
//Input[473]=8482657.07403533;
//Input[474]=8536060.61118973;
//Input[475]=8589464.14834414;
//Input[476]=8642867.68549855;
//Input[477]=8696271.22265296;
//Input[478]=8749674.75980737;
//Input[479]=8803078.29696178;
//Input[480]=8856481.83411619;
//Input[481]=8909885.3712706;
//Input[482]=8963288.90842501;
//Input[483]=9016692.44557941;
//Input[484]=9070095.98273382;
//Input[485]=9123499.51988823;
//Input[486]=9176903.05704264;
//Input[487]=9230306.59419705;
//Input[488]=9283710.13135146;
//Input[489]=9337113.66850586;
//Input[490]=9390517.20566028;
//Input[491]=9443920.74281468;
//Input[492]=9497324.27996909;
//Input[493]=9550727.8171235;
//Input[494]=9604131.35427791;
//Input[495]=9657534.89143232;
//Input[496]=9710938.42858673;
//Input[497]=9764341.96574113;
//Input[498]=9817745.50289555;
//Input[499]=9871149.04004995;
//Input[500]=9924552.57720436;
//Input[501]=9977956.11435877;
//Input[502]=10031359.6515132;
//Input[503]=10084763.1886676;
//Input[504]=10138166.725822;
//Input[505]=10191570.2629764;
//Input[506]=10244973.8001308;
//Input[507]=10298377.3372852;
//Input[508]=10351780.8744396;
//Input[509]=10405184.411594;
//Input[510]=10458587.9487485;
//Input[511]=10511991.4859029;
//Input[512]=10565395.0230573;
//Input[513]=10618798.5602117;
//Input[514]=10672202.0973661;
//Input[515]=10725605.6345205;
//Input[516]=10779009.1716749;
//Input[517]=10832412.7088293;
//Input[518]=10885816.2459837;
//Input[519]=10939219.7831381;
//Input[520]=10992623.3202925;
//Input[521]=11046026.8574469;
//Input[522]=11099430.3946014;
//Input[523]=11152833.9317558;
//Input[524]=11206237.4689102;
//Input[525]=11259641.0060646;
//Input[526]=11313044.543219;
//Input[527]=11366448.0803734;
//Input[528]=11419851.6175278;
//Input[529]=11473255.1546822;
//Input[530]=11526658.6918366;
//Input[531]=11580062.228991;
//Input[532]=11633465.7661454;
//Input[533]=11686869.3032998;
//Input[534]=11740272.8404543;
//Input[535]=11793676.3776087;
//Input[536]=11847079.9147631;
//Input[537]=11900483.4519175;
//Input[538]=11953886.9890719;
//Input[539]=12007290.5262263;
//Input[540]=12060694.0633807;
//Input[541]=12114097.6005351;
//Input[542]=12167501.1376895;
//Input[543]=12220904.6748439;
//Input[544]=12274308.2119983;
//Input[545]=12327711.7491528;
//Input[546]=12381115.2863072;
//Input[547]=12434518.8234616;
//Input[548]=12487922.360616;
//Input[549]=12541325.8977704;
//Input[550]=12594729.4349248;
//Input[551]=12648132.9720792;
//Input[552]=12701536.5092336;
//Input[553]=12754940.046388;
//Input[554]=12808343.5835424;
//Input[555]=12861747.1206968;
//Input[556]=12915150.6578513;
//Input[557]=12968554.1950057;
//Input[558]=13021957.7321601;
//Input[559]=13075361.2693145;
//Input[560]=13128764.8064689;
//Input[561]=13182168.3436233;
//Input[562]=13235571.8807777;
//Input[563]=13288975.4179321;
//Input[564]=13342378.9550865;
//Input[565]=13395782.4922409;
//Input[566]=13449186.0293953;
//Input[567]=13502589.5665497;
//Input[568]=13555993.1037042;
//Input[569]=13609396.6408586;
//Input[570]=13662800.178013;
//Input[571]=13716203.7151674;
//Input[572]=13769607.2523218;
//Input[573]=13823010.7894762;
//Input[574]=13876414.3266306;
//Input[575]=13929817.863785;
//Input[576]=13983221.4009394;
//Input[577]=14036624.9380938;
//Input[578]=14090028.4752482;
//Input[579]=14143432.0124027;
//Input[580]=14196835.5495571;
//Input[581]=14250239.0867115;
//Input[582]=14303642.6238659;
//Input[583]=14357046.1610203;
//Input[584]=14410449.6981747;
//Input[585]=14463853.2353291;
//Input[586]=14517256.7724835;
//Input[587]=14570660.3096379;
//Input[588]=14624063.8467923;
//Input[589]=14677467.3839467;
//Input[590]=14730870.9211012;
//Input[591]=14784274.4582556;
//Input[592]=14837677.99541;
//Input[593]=14891081.5325644;
//Input[594]=14944485.0697188;
//Input[595]=14997888.6068732;
//Input[596]=15051292.1440276;
//Input[597]=15104695.681182;
//Input[598]=15158099.2183364;
//Input[599]=15211502.7554908;
//Input[600]=15264906.2926452;
//Input[601]=15318309.8297996;
//Input[602]=15371713.3669541;
//Input[603]=15425116.9041085;
//Input[604]=15478520.4412629;
//Input[605]=15531923.9784173;
//Input[606]=15585327.5155717;
//Input[607]=15638731.0527261;
//Input[608]=15692134.5898805;
//Input[609]=15745538.1270349;
//Input[610]=15798941.6641893;
//Input[611]=15852345.2013437;
//Input[612]=15905748.7384981;
//Input[613]=15959152.2756525;
//Input[614]=16012555.812807;
//Input[615]=16065959.3499614;
//Input[616]=16119362.8871158;
//Input[617]=16172766.4242702;
//Input[618]=16226169.9614246;
//Input[619]=16279573.498579;
//Input[620]=16332977.0357334;
//Input[621]=16386380.5728878;
//Input[622]=16439784.1100422;
//Input[623]=16493187.6471966;
//Input[624]=16546591.184351;
//Input[625]=16599994.7215055;
//Input[626]=16653398.2586599;
//Input[627]=16706801.7958143;
//Input[628]=16760205.3329687;
//Input[629]=-16740823.1298769;

/////////////////////////////////////////////////////////////////////////
// Sin Signal
Input[0]<=0;
Input[1]<=167769;
Input[2]<=335521;
Input[3]<=503240;
Input[4]<=670909;
Input[5]<=838511;
Input[6]<=1006029;
Input[7]<=1173446;
Input[8]<=1340746;
Input[9]<=1507911;
Input[10]<=1674926;
Input[11]<=1841774;
Input[12]<=2008437;
Input[13]<=2174900;
Input[14]<=2341144;
Input[15]<=2507155;
Input[16]<=2672915;
Input[17]<=2838408;
Input[18]<=3003617;
Input[19]<=3168526;
Input[20]<=3333118;
Input[21]<=3497376;
Input[22]<=3661285;
Input[23]<=3824828;
Input[24]<=3987988;
Input[25]<=4150749;
Input[26]<=4313095;
Input[27]<=4475010;
Input[28]<=4636478;
Input[29]<=4797482;
Input[30]<=4958006;
Input[31]<=5118034;
Input[32]<=5277551;
Input[33]<=5436539;
Input[34]<=5594984;
Input[35]<=5752870;
Input[36]<=5910180;
Input[37]<=6066900;
Input[38]<=6223012;
Input[39]<=6378503;
Input[40]<=6533355;
Input[41]<=6687554;
Input[42]<=6841085;
Input[43]<=6993931;
Input[44]<=7146078;
Input[45]<=7297510;
Input[46]<=7448213;
Input[47]<=7598171;
Input[48]<=7747368;
Input[49]<=7895792;
Input[50]<=8043425;
Input[51]<=8190255;
Input[52]<=8336265;
Input[53]<=8481442;
Input[54]<=8625770;
Input[55]<=8769236;
Input[56]<=8911825;
Input[57]<=9053523;
Input[58]<=9194315;
Input[59]<=9334189;
Input[60]<=9473128;
Input[61]<=9611121;
Input[62]<=9748152;
Input[63]<=9884208;
Input[64]<=10019276;
Input[65]<=10153343;
Input[66]<=10286393;
Input[67]<=10418416;
Input[68]<=10549396;
Input[69]<=10679321;
Input[70]<=10808179;
Input[71]<=10935955;
Input[72]<=11062639;
Input[73]<=11188215;
Input[74]<=11312673;
Input[75]<=11436000;
Input[76]<=11558183;
Input[77]<=11679211;
Input[78]<=11799070;
Input[79]<=11917750;
Input[80]<=12035238;
Input[81]<=12151522;
Input[82]<=12266591;
Input[83]<=12380434;
Input[84]<=12493038;
Input[85]<=12604393;
Input[86]<=12714488;
Input[87]<=12823311;
Input[88]<=12930852;
Input[89]<=13037100;
Input[90]<=13142044;
Input[91]<=13245674;
Input[92]<=13347980;
Input[93]<=13448950;
Input[94]<=13548576;
Input[95]<=13646847;
Input[96]<=13743753;
Input[97]<=13839285;
Input[98]<=13933433;
Input[99]<=14026188;
Input[100]<=14117540;
Input[101]<=14207480;
Input[102]<=14296000;
Input[103]<=14383090;
Input[104]<=14468741;
Input[105]<=14552946;
Input[106]<=14635696;
Input[107]<=14716982;
Input[108]<=14796796;
Input[109]<=14875131;
Input[110]<=14951978;
Input[111]<=15027330;
Input[112]<=15101179;
Input[113]<=15173518;
Input[114]<=15244340;
Input[115]<=15313637;
Input[116]<=15381403;
Input[117]<=15447631;
Input[118]<=15512314;
Input[119]<=15575446;
Input[120]<=15637021;
Input[121]<=15697031;
Input[122]<=15755472;
Input[123]<=15812338;
Input[124]<=15867622;
Input[125]<=15921319;
Input[126]<=15973425;
Input[127]<=16023933;
Input[128]<=16072839;
Input[129]<=16120137;
Input[130]<=16165823;
Input[131]<=16209893;
Input[132]<=16252342;
Input[133]<=16293166;
Input[134]<=16332360;
Input[135]<=16369921;
Input[136]<=16405845;
Input[137]<=16440129;
Input[138]<=16472768;
Input[139]<=16503761;
Input[140]<=16533102;
Input[141]<=16560791;
Input[142]<=16586824;
Input[143]<=16611198;
Input[144]<=16633910;
Input[145]<=16654960;
Input[146]<=16674344;
Input[147]<=16692060;
Input[148]<=16708108;
Input[149]<=16722484;
Input[150]<=16735188;
Input[151]<=16746219;
Input[152]<=16755575;
Input[153]<=16763256;
Input[154]<=16769260;
Input[155]<=16773588;
Input[156]<=16776238;
Input[157]<=16777210;
Input[158]<=16776505;
Input[159]<=16774122;
Input[160]<=16770062;
Input[161]<=16764324;
Input[162]<=16756911;
Input[163]<=16747821;
Input[164]<=16737057;
Input[165]<=16724619;
Input[166]<=16710509;
Input[167]<=16694728;
Input[168]<=16677277;
Input[169]<=16658159;
Input[170]<=16637374;
Input[171]<=16614926;
Input[172]<=16590817;
Input[173]<=16565048;
Input[174]<=16537623;
Input[175]<=16508544;
Input[176]<=16477815;
Input[177]<=16445437;
Input[178]<=16411415;
Input[179]<=16375752;
Input[180]<=16338452;
Input[181]<=16299517;
Input[182]<=16258953;
Input[183]<=16216762;
Input[184]<=16172950;
Input[185]<=16127521;
Input[186]<=16080479;
Input[187]<=16031829;
Input[188]<=15981576;
Input[189]<=15929725;
Input[190]<=15876280;
Input[191]<=15821249;
Input[192]<=15764635;
Input[193]<=15706444;
Input[194]<=15646683;
Input[195]<=15585357;
Input[196]<=15522473;
Input[197]<=15458037;
Input[198]<=15392054;
Input[199]<=15324533;
Input[200]<=15255479;
Input[201]<=15184899;
Input[202]<=15112801;
Input[203]<=15039192;
Input[204]<=14964079;
Input[205]<=14887470;
Input[206]<=14809371;
Input[207]<=14729792;
Input[208]<=14648740;
Input[209]<=14566223;
Input[210]<=14482249;
Input[211]<=14396828;
Input[212]<=14309966;
Input[213]<=14221674;
Input[214]<=14131959;
Input[215]<=14040831;
Input[216]<=13948299;
Input[217]<=13854373;
Input[218]<=13759061;
Input[219]<=13662373;
Input[220]<=13564318;
Input[221]<=13464908;
Input[222]<=13364150;
Input[223]<=13262057;
Input[224]<=13158637;
Input[225]<=13053902;
Input[226]<=12947861;
Input[227]<=12840525;
Input[228]<=12731905;
Input[229]<=12622012;
Input[230]<=12510857;
Input[231]<=12398451;
Input[232]<=12284805;
Input[233]<=12169930;
Input[234]<=12053839;
Input[235]<=11936542;
Input[236]<=11818051;
Input[237]<=11698379;
Input[238]<=11577537;
Input[239]<=11455537;
Input[240]<=11332391;
Input[241]<=11208112;
Input[242]<=11082713;
Input[243]<=10956205;
Input[244]<=10828602;
Input[245]<=10699916;
Input[246]<=10570159;
Input[247]<=10439346;
Input[248]<=10307489;
Input[249]<=10174601;
Input[250]<=10040696;
Input[251]<=9905787;
Input[252]<=9769887;
Input[253]<=9633010;
Input[254]<=9495169;
Input[255]<=9356380;
Input[256]<=9216654;
Input[257]<=9076007;
Input[258]<=8934453;
Input[259]<=8792005;
Input[260]<=8648677;
Input[261]<=8504485;
Input[262]<=8359443;
Input[263]<=8213564;
Input[264]<=8066864;
Input[265]<=7919358;
Input[266]<=7771059;
Input[267]<=7621984;
Input[268]<=7472146;
Input[269]<=7321561;
Input[270]<=7170244;
Input[271]<=7018210;
Input[272]<=6865474;
Input[273]<=6712052;
Input[274]<=6557958;
Input[275]<=6403208;
Input[276]<=6247819;
Input[277]<=6091804;
Input[278]<=5935180;
Input[279]<=5777963;
Input[280]<=5620168;
Input[281]<=5461811;
Input[282]<=5302908;
Input[283]<=5143474;
Input[284]<=4983526;
Input[285]<=4823080;
Input[286]<=4662152;
Input[287]<=4500757;
Input[288]<=4338912;
Input[289]<=4176634;
Input[290]<=4013937;
Input[291]<=3850839;
Input[292]<=3687357;
Input[293]<=3523505;
Input[294]<=3359301;
Input[295]<=3194761;
Input[296]<=3029902;
Input[297]<=2864740;
Input[298]<=2699291;
Input[299]<=2533572;
Input[300]<=2367600;
Input[301]<=2201392;
Input[302]<=2034963;
Input[303]<=1868330;
Input[304]<=1701511;
Input[305]<=1534522;
Input[306]<=1367379;
Input[307]<=1200099;
Input[308]<=1032700;
Input[309]<=865197;
Input[310]<=697607;
Input[311]<=529948;
Input[312]<=362236;
Input[313]<=194488;
Input[314]<=26720;
Input[315]<=-141050;
Input[316]<=-308806;
Input[317]<=-476532;
Input[318]<=-644209;
Input[319]<=-811823;
Input[320]<=-979355;
Input[321]<=-1146789;
Input[322]<=-1314109;
Input[323]<=-1481297;
Input[324]<=-1648337;
Input[325]<=-1815213;
Input[326]<=-1981906;
Input[327]<=-2148402;
Input[328]<=-2314683;
Input[329]<=-2480732;
Input[330]<=-2646533;
Input[331]<=-2812070;
Input[332]<=-2977325;
Input[333]<=-3142283;
Input[334]<=-3306926;
Input[335]<=-3471239;
Input[336]<=-3635204;
Input[337]<=-3798806;
Input[338]<=-3962028;
Input[339]<=-4124854;
Input[340]<=-4287268;
Input[341]<=-4449253;
Input[342]<=-4610792;
Input[343]<=-4771871;
Input[344]<=-4932473;
Input[345]<=-5092581;
Input[346]<=-5252180;
Input[347]<=-5411254;
Input[348]<=-5569787;
Input[349]<=-5727762;
Input[350]<=-5885165;
Input[351]<=-6041980;
Input[352]<=-6198190;
Input[353]<=-6353781;
Input[354]<=-6508736;
Input[355]<=-6663040;
Input[356]<=-6816678;
Input[357]<=-6969634;
Input[358]<=-7121894;
Input[359]<=-7273441;
Input[360]<=-7424261;
Input[361]<=-7574338;
Input[362]<=-7723658;
Input[363]<=-7872205;
Input[364]<=-8019966;
Input[365]<=-8166924;
Input[366]<=-8313066;
Input[367]<=-8458376;
Input[368]<=-8602841;
Input[369]<=-8746445;
Input[370]<=-8889175;
Input[371]<=-9031016;
Input[372]<=-9171953;
Input[373]<=-9311974;
Input[374]<=-9451063;
Input[375]<=-9589207;
Input[376]<=-9726392;
Input[377]<=-9862605;
Input[378]<=-9997831;
Input[379]<=-10132058;
Input[380]<=-10265271;
Input[381]<=-10397458;
Input[382]<=-10528606;
Input[383]<=-10658700;
Input[384]<=-10787728;
Input[385]<=-10915678;
Input[386]<=-11042536;
Input[387]<=-11168290;
Input[388]<=-11292927;
Input[389]<=-11416435;
Input[390]<=-11538801;
Input[391]<=-11660013;
Input[392]<=-11780059;
Input[393]<=-11898928;
Input[394]<=-12016606;
Input[395]<=-12133083;
Input[396]<=-12248346;
Input[397]<=-12362385;
Input[398]<=-12475187;
Input[399]<=-12586742;
Input[400]<=-12697038;
Input[401]<=-12806065;
Input[402]<=-12913811;
Input[403]<=-13020265;
Input[404]<=-13125418;
Input[405]<=-13229258;
Input[406]<=-13331775;
Input[407]<=-13432959;
Input[408]<=-13532800;
Input[409]<=-13631287;
Input[410]<=-13728411;
Input[411]<=-13824163;
Input[412]<=-13918532;
Input[413]<=-14011509;
Input[414]<=-14103085;
Input[415]<=-14193251;
Input[416]<=-14281997;
Input[417]<=-14369315;
Input[418]<=-14455197;
Input[419]<=-14539633;
Input[420]<=-14622614;
Input[421]<=-14704134;
Input[422]<=-14784183;
Input[423]<=-14862754;
Input[424]<=-14939839;
Input[425]<=-15015429;
Input[426]<=-15089518;
Input[427]<=-15162098;
Input[428]<=-15233162;
Input[429]<=-15302703;
Input[430]<=-15370713;
Input[431]<=-15437187;
Input[432]<=-15502116;
Input[433]<=-15565496;
Input[434]<=-15627318;
Input[435]<=-15687579;
Input[436]<=-15746270;
Input[437]<=-15803387;
Input[438]<=-15858923;
Input[439]<=-15912874;
Input[440]<=-15965233;
Input[441]<=-16015996;
Input[442]<=-16065157;
Input[443]<=-16112712;
Input[444]<=-16158655;
Input[445]<=-16202983;
Input[446]<=-16245690;
Input[447]<=-16286773;
Input[448]<=-16326227;
Input[449]<=-16364048;
Input[450]<=-16400233;
Input[451]<=-16434779;
Input[452]<=-16467680;
Input[453]<=-16498935;
Input[454]<=-16528540;
Input[455]<=-16556492;
Input[456]<=-16582789;
Input[457]<=-16607427;
Input[458]<=-16630404;
Input[459]<=-16651719;
Input[460]<=-16671368;
Input[461]<=-16689350;
Input[462]<=-16705664;
Input[463]<=-16720306;
Input[464]<=-16733277;
Input[465]<=-16744574;
Input[466]<=-16754197;
Input[467]<=-16762145;
Input[468]<=-16768416;
Input[469]<=-16773011;
Input[470]<=-16775928;
Input[471]<=-16777168;
Input[472]<=-16776730;
Input[473]<=-16774614;
Input[474]<=-16770821;
Input[475]<=-16765350;
Input[476]<=-16758204;
Input[477]<=-16749381;
Input[478]<=-16738884;
Input[479]<=-16726712;
Input[480]<=-16712868;
Input[481]<=-16697353;
Input[482]<=-16680168;
Input[483]<=-16661315;
Input[484]<=-16640796;
Input[485]<=-16618613;
Input[486]<=-16594768;
Input[487]<=-16569263;
Input[488]<=-16542102;
Input[489]<=-16513286;
Input[490]<=-16482819;
Input[491]<=-16450704;
Input[492]<=-16416944;
Input[493]<=-16381542;
Input[494]<=-16344502;
Input[495]<=-16305827;
Input[496]<=-16265522;
Input[497]<=-16223591;
Input[498]<=-16180037;
Input[499]<=-16134865;
Input[500]<=-16088079;
Input[501]<=-16039685;
Input[502]<=-15989687;
Input[503]<=-15938090;
Input[504]<=-15884899;
Input[505]<=-15830119;
Input[506]<=-15773757;
Input[507]<=-15715817;
Input[508]<=-15656306;
Input[509]<=-15595229;
Input[510]<=-15532592;
Input[511]<=-15468403;
Input[512]<=-15402666;
Input[513]<=-15335389;
Input[514]<=-15266579;
Input[515]<=-15196242;
Input[516]<=-15124386;
Input[517]<=-15051017;
Input[518]<=-14976142;
Input[519]<=-14899771;
Input[520]<=-14821909;
Input[521]<=-14742565;
Input[522]<=-14661747;
Input[523]<=-14579463;
Input[524]<=-14495721;
Input[525]<=-14410529;
Input[526]<=-14323896;
Input[527]<=-14235831;
Input[528]<=-14146342;
Input[529]<=-14055439;
Input[530]<=-13963130;
Input[531]<=-13869425;
Input[532]<=-13774333;
Input[533]<=-13677863;
Input[534]<=-13580026;
Input[535]<=-13480831;
Input[536]<=-13380287;
Input[537]<=-13278406;
Input[538]<=-13175197;
Input[539]<=-13070670;
Input[540]<=-12964836;
Input[541]<=-12857706;
Input[542]<=-12749290;
Input[543]<=-12639599;
Input[544]<=-12528644;
Input[545]<=-12416436;
Input[546]<=-12302987;
Input[547]<=-12188307;
Input[548]<=-12072409;
Input[549]<=-11955303;
Input[550]<=-11837002;
Input[551]<=-11717517;
Input[552]<=-11596860;
Input[553]<=-11475044;
Input[554]<=-11352080;
Input[555]<=-11227981;
Input[556]<=-11102759;
Input[557]<=-10976427;
Input[558]<=-10848998;
Input[559]<=-10720483;
Input[560]<=-10590896;
Input[561]<=-10460251;
Input[562]<=-10328559;
Input[563]<=-10195834;
Input[564]<=-10062090;
Input[565]<=-9927340;
Input[566]<=-9791597;
Input[567]<=-9654874;
Input[568]<=-9517187;
Input[569]<=-9378547;
Input[570]<=-9238970;
Input[571]<=-9098469;
Input[572]<=-8957058;
Input[573]<=-8814751;
Input[574]<=-8671563;
Input[575]<=-8527507;
Input[576]<=-8382599;
Input[577]<=-8236853;
Input[578]<=-8090283;
Input[579]<=-7942904;
Input[580]<=-7794731;
Input[581]<=-7645778;
Input[582]<=-7496060;
Input[583]<=-7345594;
Input[584]<=-7194392;
Input[585]<=-7042471;
Input[586]<=-6889846;
Input[587]<=-6736532;
Input[588]<=-6582544;
Input[589]<=-6427898;
Input[590]<=-6272609;
Input[591]<=-6116693;
Input[592]<=-5960165;
Input[593]<=-5803041;
Input[594]<=-5645337;
Input[595]<=-5487069;
Input[596]<=-5328251;
Input[597]<=-5168901;
Input[598]<=-5009034;
Input[599]<=-4848666;
Input[600]<=-4687814;
Input[601]<=-4526492;
Input[602]<=-4364718;
Input[603]<=-4202507;
Input[604]<=-4039876;
Input[605]<=-3876841;
Input[606]<=-3713419;
Input[607]<=-3549625;
Input[608]<=-3385476;
Input[609]<=-3220989;
Input[610]<=-3056179;
Input[611]<=-2891064;
Input[612]<=-2725660;
Input[613]<=-2559983;
Input[614]<=-2394050;
Input[615]<=-2227878;
Input[616]<=-2061483;
Input[617]<=-1894882;
Input[618]<=-1728091;
Input[619]<=-1561128;
Input[620]<=-1394008;
Input[621]<=-1226749;
Input[622]<=-1059368;
Input[623]<=-891880;
Input[624]<=-724304;
Input[625]<=-556654;
Input[626]<=-388950;
Input[627]<=-221206;
Input[628]<=-53440;
Input[629]<=114330;
Input[630]<=282090;
Input[631]<=449821;
Input[632]<=617508;
Input[633]<=785133;
Input[634]<=952679;
Input[635]<=1120130;
Input[636]<=1287469;
Input[637]<=1454679;
Input[638]<=1621744;
Input[639]<=1788647;
Input[640]<=1955371;
Input[641]<=2121899;
Input[642]<=2288215;
Input[643]<=2454302;
Input[644]<=2620144;
Input[645]<=2785724;
Input[646]<=2951025;
Input[647]<=3116031;
Input[648]<=3280726;
Input[649]<=3445092;
Input[650]<=3609114;
Input[651]<=3772775;
Input[652]<=3936059;
Input[653]<=4098949;
Input[654]<=4261429;
Input[655]<=4423483;
Input[656]<=4585095;
Input[657]<=4746248;
Input[658]<=4906927;
Input[659]<=5067115;
Input[660]<=5226796;
Input[661]<=5385955;
Input[662]<=5544575;
Input[663]<=5702640;
Input[664]<=5860136;
Input[665]<=6017045;
Input[666]<=6173352;
Input[667]<=6329043;
Input[668]<=6484100;
Input[669]<=6638509;
Input[670]<=6792254;
Input[671]<=6945320;
Input[672]<=7097691;
Input[673]<=7249353;
Input[674]<=7400290;
Input[675]<=7550486;
Input[676]<=7699928;
Input[677]<=7848599;
Input[678]<=7996486;
Input[679]<=8143573;
Input[680]<=8289846;
Input[681]<=8435290;
Input[682]<=8579890;
Input[683]<=8723632;
Input[684]<=8866502;
Input[685]<=9008485;
Input[686]<=9149568;
Input[687]<=9289735;
Input[688]<=9428974;
Input[689]<=9567269;
Input[690]<=9704608;
Input[691]<=9840977;
Input[692]<=9976361;
Input[693]<=10110748;
Input[694]<=10244124;
Input[695]<=10376475;
Input[696]<=10507788;
Input[697]<=10638051;
Input[698]<=10767250;
Input[699]<=10895373;
Input[700]<=11022406;
Input[701]<=11148336;
Input[702]<=11273152;
Input[703]<=11396840;
Input[704]<=11519389;
Input[705]<=11640786;
Input[706]<=11761019;
Input[707]<=11880075;
Input[708]<=11997944;
Input[709]<=12114613;
Input[710]<=12230071;
Input[711]<=12344305;
Input[712]<=12457305;
Input[713]<=12569059;
Input[714]<=12679557;
Input[715]<=12788786;
Input[716]<=12896737;
Input[717]<=13003398;
Input[718]<=13108758;
Input[719]<=13212808;
Input[720]<=13315537;
Input[721]<=13416934;
Input[722]<=13516989;
Input[723]<=13615692;
Input[724]<=13713034;
Input[725]<=13809005;
Input[726]<=13903595;
Input[727]<=13996795;
Input[728]<=14088594;
Input[729]<=14178985;
Input[730]<=14267958;
Input[731]<=14355505;
Input[732]<=14441615;
Input[733]<=14526282;
Input[734]<=14609496;
Input[735]<=14691249;
Input[736]<=14771533;
Input[737]<=14850340;
Input[738]<=14927662;
Input[739]<=15003491;
Input[740]<=15077819;
Input[741]<=15150640;
Input[742]<=15221946;
Input[743]<=15291730;
Input[744]<=15359984;
Input[745]<=15426703;
Input[746]<=15491879;
Input[747]<=15555505;
Input[748]<=15617577;
Input[749]<=15678086;
Input[750]<=15737028;
Input[751]<=15794396;
Input[752]<=15850184;
Input[753]<=15904388;
Input[754]<=15957001;
Input[755]<=16008018;
Input[756]<=16057435;
Input[757]<=16105246;
Input[758]<=16151446;
Input[759]<=16196031;
Input[760]<=16238997;
Input[761]<=16280339;
Input[762]<=16320052;
Input[763]<=16358134;
Input[764]<=16394580;
Input[765]<=16429387;
Input[766]<=16462550;
Input[767]<=16494068;
Input[768]<=16523935;
Input[769]<=16552151;
Input[770]<=16578711;
Input[771]<=16603614;
Input[772]<=16626856;
Input[773]<=16648436;
Input[774]<=16668350;
Input[775]<=16686598;
Input[776]<=16703177;
Input[777]<=16718086;
Input[778]<=16731323;
Input[779]<=16742887;
Input[780]<=16752777;
Input[781]<=16760991;
Input[782]<=16767530;
Input[783]<=16772391;
Input[784]<=16775576;
Input[785]<=16777083;
Input[786]<=16776912;
Input[787]<=16775063;
Input[788]<=16771537;
Input[789]<=16766334;
Input[790]<=16759454;
Input[791]<=16750898;
Input[792]<=16740668;
Input[793]<=16728763;
Input[794]<=16715185;
Input[795]<=16699936;
Input[796]<=16683017;
Input[797]<=16664429;
Input[798]<=16644175;
Input[799]<=16622257;
Input[800]<=16598677;
Input[801]<=16573436;
Input[802]<=16546538;
Input[803]<=16517986;
Input[804]<=16487782;
Input[805]<=16455929;
Input[806]<=16422431;
Input[807]<=16387290;
Input[808]<=16350510;
Input[809]<=16312096;
Input[810]<=16272050;
Input[811]<=16230378;
Input[812]<=16187082;
Input[813]<=16142167;
Input[814]<=16095638;
Input[815]<=16047500;
Input[816]<=15997757;
Input[817]<=15946414;
Input[818]<=15893477;
Input[819]<=15838950;
Input[820]<=15782839;
Input[821]<=15725150;
Input[822]<=15665889;
Input[823]<=15605061;
Input[824]<=15542672;
Input[825]<=15478730;
Input[826]<=15413239;
Input[827]<=15346207;
Input[828]<=15277641;
Input[829]<=15207546;
Input[830]<=15135931;
Input[831]<=15062803;
Input[832]<=14988168;
Input[833]<=14912034;
Input[834]<=14834409;
Input[835]<=14755301;
Input[836]<=14674717;
Input[837]<=14592666;
Input[838]<=14509155;
Input[839]<=14424194;
Input[840]<=14337790;
Input[841]<=14249952;
Input[842]<=14160690;
Input[843]<=14070011;
Input[844]<=13977925;
Input[845]<=13884442;
Input[846]<=13789570;
Input[847]<=13693319;
Input[848]<=13595699;
Input[849]<=13496720;
Input[850]<=13396390;
Input[851]<=13294721;
Input[852]<=13191723;
Input[853]<=13087405;
Input[854]<=12981779;
Input[855]<=12874854;
Input[856]<=12766643;
Input[857]<=12657154;
Input[858]<=12546400;
Input[859]<=12434391;
Input[860]<=12321138;
Input[861]<=12206654;
Input[862]<=12090949;
Input[863]<=11974034;
Input[864]<=11855923;
Input[865]<=11736626;
Input[866]<=11616155;
Input[867]<=11494522;
Input[868]<=11371740;
Input[869]<=11247821;
Input[870]<=11122777;
Input[871]<=10996621;
Input[872]<=10869366;
Input[873]<=10741023;
Input[874]<=10611606;
Input[875]<=10481128;
Input[876]<=10349602;
Input[877]<=10217041;
Input[878]<=10083459;
Input[879]<=9948867;
Input[880]<=9813282;
Input[881]<=9676714;
Input[882]<=9539179;
Input[883]<=9400691;
Input[884]<=9261262;
Input[885]<=9120907;
Input[886]<=8979640;
Input[887]<=8837475;
Input[888]<=8694426;
Input[889]<=8550508;
Input[890]<=8405735;
Input[891]<=8260121;
Input[892]<=8113681;
Input[893]<=7966430;
Input[894]<=7818382;
Input[895]<=7669552;
Input[896]<=7519956;
Input[897]<=7369607;
Input[898]<=7218522;
Input[899]<=7066714;
Input[900]<=6914200;
Input[901]<=6760995;
Input[902]<=6607113;
Input[903]<=6452571;
Input[904]<=6297384;
Input[905]<=6141566;
Input[906]<=5985135;
Input[907]<=5828105;
Input[908]<=5670492;
Input[909]<=5512313;
Input[910]<=5353582;
Input[911]<=5194315;
Input[912]<=5034530;
Input[913]<=4874240;
Input[914]<=4713464;
Input[915]<=4552216;
Input[916]<=4390513;
Input[917]<=4228370;
Input[918]<=4065805;
Input[919]<=3902834;
Input[920]<=3739472;
Input[921]<=3575736;
Input[922]<=3411642;
Input[923]<=3247208;
Input[924]<=3082449;
Input[925]<=2917381;
Input[926]<=2752022;
Input[927]<=2586387;
Input[928]<=2420494;
Input[929]<=2254359;
Input[930]<=2087998;
Input[931]<=1921429;
Input[932]<=1754667;
Input[933]<=1587730;
Input[934]<=1420634;
Input[935]<=1253397;
Input[936]<=1086033;
Input[937]<=918562;
Input[938]<=750998;
Input[939]<=583359;
Input[940]<=415662;
Input[941]<=247924;
Input[942]<=80160;
Input[943]<=-87610;
Input[944]<=-255373;
Input[945]<=-423110;
Input[946]<=-590805;
Input[947]<=-758441;
Input[948]<=-926001;
Input[949]<=-1093468;
Input[950]<=-1260826;
Input[951]<=-1428058;
Input[952]<=-1595147;
Input[953]<=-1762077;
Input[954]<=-1928830;
Input[955]<=-2095391;
Input[956]<=-2261741;
Input[957]<=-2427866;
Input[958]<=-2593748;
Input[959]<=-2759371;
Input[960]<=-2924718;
Input[961]<=-3089772;
Input[962]<=-3254517;
Input[963]<=-3418937;
Input[964]<=-3583015;
Input[965]<=-3746734;
Input[966]<=-3910079;
Input[967]<=-4073033;
Input[968]<=-4235580;
Input[969]<=-4397703;
Input[970]<=-4559386;
Input[971]<=-4720614;
Input[972]<=-4881369;
Input[973]<=-5041636;
Input[974]<=-5201399;
Input[975]<=-5360642;
Input[976]<=-5519349;
Input[977]<=-5677504;
Input[978]<=-5835091;
Input[979]<=-5992095;
Input[980]<=-6148499;
Input[981]<=-6304289;
Input[982]<=-6459448;
Input[983]<=-6613961;
Input[984]<=-6767813;
Input[985]<=-6920988;
Input[986]<=-7073471;
Input[987]<=-7225247;
Input[988]<=-7376300;
Input[989]<=-7526615;
Input[990]<=-7676178;
Input[991]<=-7824973;
Input[992]<=-7972986;
Input[993]<=-8120201;
Input[994]<=-8266605;
Input[995]<=-8412182;
Input[996]<=-8556917;
Input[997]<=-8700797;
Input[998]<=-8843807;
Input[999]<=-8985932;
Input[1000]<=-9127159;
Input[1001]<=-9267473;
Input[1002]<=-9406861;
Input[1003]<=-9545307;
Input[1004]<=-9682800;
Input[1005]<=-9819324;
Input[1006]<=-9954866;
Input[1007]<=-10089412;
Input[1008]<=-10222950;
Input[1009]<=-10355465;
Input[1010]<=-10486945;
Input[1011]<=-10617376;
Input[1012]<=-10746745;
Input[1013]<=-10875040;
Input[1014]<=-11002247;
Input[1015]<=-11128354;
Input[1016]<=-11253348;
Input[1017]<=-11377217;
Input[1018]<=-11499948;
Input[1019]<=-11621529;
Input[1020]<=-11741948;
Input[1021]<=-11861193;
Input[1022]<=-11979252;
Input[1023]<=-12096113;
Input[1024]<=-12211764;
Input[1025]<=-12326194;
Input[1026]<=-12439391;
Input[1027]<=-12551345;
Input[1028]<=-12662043;
Input[1029]<=-12771475;
Input[1030]<=-12879630;
Input[1031]<=-12986497;
Input[1032]<=-13092066;
Input[1033]<=-13196325;
Input[1034]<=-13299264;
Input[1035]<=-13400874;
Input[1036]<=-13501144;
Input[1037]<=-13600063;
Input[1038]<=-13697623;
Input[1039]<=-13793813;
Input[1040]<=-13888623;
Input[1041]<=-13982045;
Input[1042]<=-14074068;
Input[1043]<=-14164684;
Input[1044]<=-14253883;
Input[1045]<=-14341657;
Input[1046]<=-14427997;
Input[1047]<=-14512895;
Input[1048]<=-14596341;
Input[1049]<=-14678327;
Input[1050]<=-14758845;
Input[1051]<=-14837888;
Input[1052]<=-14915447;
Input[1053]<=-14991514;
Input[1054]<=-15066082;
Input[1055]<=-15139144;
Input[1056]<=-15210691;
Input[1057]<=-15280718;
Input[1058]<=-15349216;
Input[1059]<=-15416180;
Input[1060]<=-15481602;
Input[1061]<=-15545476;
Input[1062]<=-15607795;
Input[1063]<=-15668554;
Input[1064]<=-15727746;
Input[1065]<=-15785365;
Input[1066]<=-15841405;
Input[1067]<=-15895861;
Input[1068]<=-15948728;
Input[1069]<=-16000000;
Input[1070]<=-16049672;
Input[1071]<=-16097739;
Input[1072]<=-16144196;
Input[1073]<=-16189039;
Input[1074]<=-16232263;
Input[1075]<=-16273863;
Input[1076]<=-16313837;
Input[1077]<=-16352178;
Input[1078]<=-16388885;
Input[1079]<=-16423953;
Input[1080]<=-16457379;
Input[1081]<=-16489158;
Input[1082]<=-16519289;
Input[1083]<=-16547768;
Input[1084]<=-16574592;
Input[1085]<=-16599759;
Input[1086]<=-16623266;
Input[1087]<=-16645110;
Input[1088]<=-16665290;
Input[1089]<=-16683803;
Input[1090]<=-16700649;
Input[1091]<=-16715824;
Input[1092]<=-16729327;
Input[1093]<=-16741158;
Input[1094]<=-16751314;
Input[1095]<=-16759795;
Input[1096]<=-16766601;
Input[1097]<=-16771729;
Input[1098]<=-16775181;
Input[1099]<=-16776955;
Input[1100]<=-16777051;
Input[1101]<=-16775470;
Input[1102]<=-16772211;
Input[1103]<=-16767275;
Input[1104]<=-16760662;
Input[1105]<=-16752373;
Input[1106]<=-16742409;
Input[1107]<=-16730771;
Input[1108]<=-16717460;
Input[1109]<=-16702476;
Input[1110]<=-16685823;
Input[1111]<=-16667501;
Input[1112]<=-16647513;
Input[1113]<=-16625859;
Input[1114]<=-16602543;
Input[1115]<=-16577567;
Input[1116]<=-16550933;
Input[1117]<=-16522644;
Input[1118]<=-16492703;
Input[1119]<=-16461112;
Input[1120]<=-16427876;
Input[1121]<=-16392996;
Input[1122]<=-16356478;
Input[1123]<=-16318323;
Input[1124]<=-16278537;
Input[1125]<=-16237123;
Input[1126]<=-16194086;
Input[1127]<=-16149429;
Input[1128]<=-16103157;
Input[1129]<=-16055274;
Input[1130]<=-16005787;
Input[1131]<=-15954698;
Input[1132]<=-15902014;
Input[1133]<=-15847740;
Input[1134]<=-15791882;
Input[1135]<=-15734444;
Input[1136]<=-15675432;
Input[1137]<=-15614853;
Input[1138]<=-15552713;
Input[1139]<=-15489017;
Input[1140]<=-15423773;
Input[1141]<=-15356986;
Input[1142]<=-15288663;
Input[1143]<=-15218812;
Input[1144]<=-15147439;
Input[1145]<=-15074551;
Input[1146]<=-15000155;
Input[1147]<=-14924260;
Input[1148]<=-14846872;
Input[1149]<=-14767999;
Input[1150]<=-14687650;
Input[1151]<=-14605832;
Input[1152]<=-14522553;
Input[1153]<=-14437822;
Input[1154]<=-14351647;
Input[1155]<=-14264037;
Input[1156]<=-14175001;
Input[1157]<=-14084548;
Input[1158]<=-13992685;
Input[1159]<=-13899424;
Input[1160]<=-13804773;
Input[1161]<=-13708741;
Input[1162]<=-13611338;
Input[1163]<=-13512574;
Input[1164]<=-13412459;
Input[1165]<=-13311003;
Input[1166]<=-13208216;
Input[1167]<=-13104107;
Input[1168]<=-12998689;
Input[1169]<=-12891970;
Input[1170]<=-12783963;
Input[1171]<=-12674677;
Input[1172]<=-12564123;
Input[1173]<=-12452313;
Input[1174]<=-12339258;
Input[1175]<=-12224969;
Input[1176]<=-12109458;
Input[1177]<=-11992735;
Input[1178]<=-11874814;
Input[1179]<=-11755704;
Input[1180]<=-11635420;
Input[1181]<=-11513971;
Input[1182]<=-11391372;
Input[1183]<=-11267633;
Input[1184]<=-11142767;
Input[1185]<=-11016788;
Input[1186]<=-10889706;
Input[1187]<=-10761536;
Input[1188]<=-10632289;
Input[1189]<=-10501979;
Input[1190]<=-10370619;
Input[1191]<=-10238222;
Input[1192]<=-10104801;
Input[1193]<=-9970370;
Input[1194]<=-9834942;
Input[1195]<=-9698530;
Input[1196]<=-9561148;
Input[1197]<=-9422810;
Input[1198]<=-9283530;
Input[1199]<=-9143322;
Input[1200]<=-9002199;
Input[1201]<=-8860176;
Input[1202]<=-8717267;
Input[1203]<=-8573487;
Input[1204]<=-8428849;
Input[1205]<=-8283368;
Input[1206]<=-8137059;
Input[1207]<=-7989936;
Input[1208]<=-7842014;
Input[1209]<=-7693308;
Input[1210]<=-7543832;
Input[1211]<=-7393602;
Input[1212]<=-7242633;
Input[1213]<=-7090940;
Input[1214]<=-6938537;
Input[1215]<=-6785441;
Input[1216]<=-6631666;
Input[1217]<=-6477228;
Input[1218]<=-6322142;
Input[1219]<=-6166424;
Input[1220]<=-6010090;
Input[1221]<=-5853154;
Input[1222]<=-5695633;
Input[1223]<=-5537542;
Input[1224]<=-5378898;
Input[1225]<=-5219716;
Input[1226]<=-5060012;
Input[1227]<=-4899802;
Input[1228]<=-4739102;
Input[1229]<=-4577928;
Input[1230]<=-4416296;
Input[1231]<=-4254223;
Input[1232]<=-4091724;
Input[1233]<=-3928816;
Input[1234]<=-3765515;
Input[1235]<=-3601838;
Input[1236]<=-3437800;
Input[1237]<=-3273419;
Input[1238]<=-3108710;
Input[1239]<=-2943690;
Input[1240]<=-2778377;
Input[1241]<=-2612785;
Input[1242]<=-2446932;
Input[1243]<=-2280834;
Input[1244]<=-2114508;
Input[1245]<=-1947971;
Input[1246]<=-1781239;
Input[1247]<=-1614329;
Input[1248]<=-1447257;
Input[1249]<=-1280041;
Input[1250]<=-1112696;
Input[1251]<=-945241;
Input[1252]<=-777691;
Input[1253]<=-610063;
Input[1254]<=-442374;
Input[1255]<=-274641;
Input[1256]<=-106880;
Input[1257]<=60890;
Input[1258]<=228656;
Input[1259]<=396398;
Input[1260]<=564101;
Input[1261]<=731747;
Input[1262]<=899320;
Input[1263]<=1066803;
Input[1264]<=1234180;
Input[1265]<=1401433;
Input[1266]<=1568546;
Input[1267]<=1735502;
Input[1268]<=1902284;
Input[1269]<=2068877;
Input[1270]<=2235262;
Input[1271]<=2401424;
Input[1272]<=2567346;
Input[1273]<=2733011;
Input[1274]<=2898403;
Input[1275]<=3063505;
Input[1276]<=3228300;
Input[1277]<=3392773;
Input[1278]<=3556906;
Input[1279]<=3720684;
Input[1280]<=3884090;
Input[1281]<=4047107;
Input[1282]<=4209720;
Input[1283]<=4371911;
Input[1284]<=4533666;
Input[1285]<=4694967;
Input[1286]<=4855798;
Input[1287]<=5016144;
Input[1288]<=5175989;
Input[1289]<=5335316;
Input[1290]<=5494109;
Input[1291]<=5652353;
Input[1292]<=5810031;
Input[1293]<=5967129;
Input[1294]<=6123630;
Input[1295]<=6279519;
Input[1296]<=6434779;
Input[1297]<=6589396;
Input[1298]<=6743355;
Input[1299]<=6896638;
Input[1300]<=7049233;
Input[1301]<=7201122;
Input[1302]<=7352291;
Input[1303]<=7502725;
Input[1304]<=7652409;
Input[1305]<=7801327;
Input[1306]<=7949466;
Input[1307]<=8096809;
Input[1308]<=8243343;
Input[1309]<=8389052;
Input[1310]<=8533923;
Input[1311]<=8677940;
Input[1312]<=8821089;
Input[1313]<=8963356;
Input[1314]<=9104727;
Input[1315]<=9245188;
Input[1316]<=9384724;
Input[1317]<=9523321;
Input[1318]<=9660966;
Input[1319]<=9797645;
Input[1320]<=9933345;
Input[1321]<=10068051;
Input[1322]<=10201750;
Input[1323]<=10334429;
Input[1324]<=10466074;
Input[1325]<=10596673;
Input[1326]<=10726213;
Input[1327]<=10854679;
Input[1328]<=10982061;
Input[1329]<=11108344;
Input[1330]<=11233516;
Input[1331]<=11357565;
Input[1332]<=11480478;
Input[1333]<=11602243;
Input[1334]<=11722848;
Input[1335]<=11842281;
Input[1336]<=11960529;
Input[1337]<=12077581;
Input[1338]<=12193426;
Input[1339]<=12308051;
Input[1340]<=12421446;
Input[1341]<=12533598;
Input[1342]<=12644497;
Input[1343]<=12754132;
Input[1344]<=12862491;
Input[1345]<=12969564;
Input[1346]<=13075340;
Input[1347]<=13179808;
Input[1348]<=13282959;
Input[1349]<=13384781;
Input[1350]<=13485264;
Input[1351]<=13584400;
Input[1352]<=13682176;
Input[1353]<=13778585;
Input[1354]<=13873616;
Input[1355]<=13967259;
Input[1356]<=14059506;
Input[1357]<=14150346;
Input[1358]<=14239772;
Input[1359]<=14327774;
Input[1360]<=14414343;
Input[1361]<=14499470;
Input[1362]<=14583148;
Input[1363]<=14665367;
Input[1364]<=14746120;
Input[1365]<=14825398;
Input[1366]<=14903194;
Input[1367]<=14979499;
Input[1368]<=15054307;
Input[1369]<=15127609;
Input[1370]<=15199398;
Input[1371]<=15269667;
Input[1372]<=15338410;
Input[1373]<=15405618;
Input[1374]<=15471286;
Input[1375]<=15535407;
Input[1376]<=15597974;
Input[1377]<=15658982;
Input[1378]<=15718424;
Input[1379]<=15776293;
Input[1380]<=15832586;
Input[1381]<=15887295;
Input[1382]<=15940415;
Input[1383]<=15991941;
Input[1384]<=16041868;
Input[1385]<=16090191;
Input[1386]<=16136905;
Input[1387]<=16182005;
Input[1388]<=16225487;
Input[1389]<=16267347;
Input[1390]<=16307579;
Input[1391]<=16346181;
Input[1392]<=16383149;
Input[1393]<=16418478;
Input[1394]<=16452165;
Input[1395]<=16484207;
Input[1396]<=16514601;
Input[1397]<=16543343;
Input[1398]<=16570431;
Input[1399]<=16595862;
Input[1400]<=16619633;
Input[1401]<=16641742;
Input[1402]<=16662188;
Input[1403]<=16680967;
Input[1404]<=16698077;
Input[1405]<=16713519;
Input[1406]<=16727288;
Input[1407]<=16739385;
Input[1408]<=16749808;
Input[1409]<=16758557;
Input[1410]<=16765629;
Input[1411]<=16771025;
Input[1412]<=16774743;
Input[1413]<=16776785;
Input[1414]<=16777148;
Input[1415]<=16775834;
Input[1416]<=16772842;
Input[1417]<=16768173;
Input[1418]<=16761828;
Input[1419]<=16753806;
Input[1420]<=16744108;
Input[1421]<=16732737;
Input[1422]<=16719692;
Input[1423]<=16704975;
Input[1424]<=16688587;
Input[1425]<=16670531;
Input[1426]<=16650808;
Input[1427]<=16629419;
Input[1428]<=16606368;
Input[1429]<=16581656;
Input[1430]<=16555286;
Input[1431]<=16527260;
Input[1432]<=16497582;
Input[1433]<=16466254;
Input[1434]<=16433279;
Input[1435]<=16398661;
Input[1436]<=16362403;
Input[1437]<=16324509;
Input[1438]<=16284983;
Input[1439]<=16243828;
Input[1440]<=16201049;
Input[1441]<=16156649;
Input[1442]<=16110634;
Input[1443]<=16063008;
Input[1444]<=16013776;
Input[1445]<=15962942;
Input[1446]<=15910512;
Input[1447]<=15856491;
Input[1448]<=15800884;
Input[1449]<=15743697;
Input[1450]<=15684936;
Input[1451]<=15624606;
Input[1452]<=15562714;
Input[1453]<=15499266;
Input[1454]<=15434267;
Input[1455]<=15367726;
Input[1456]<=15299647;
Input[1457]<=15230039;
Input[1458]<=15158907;
Input[1459]<=15086260;
Input[1460]<=15012104;
Input[1461]<=14936447;
Input[1462]<=14859296;
Input[1463]<=14780660;
Input[1464]<=14700545;
Input[1465]<=14618960;
Input[1466]<=14535914;
Input[1467]<=14451414;
Input[1468]<=14365468;
Input[1469]<=14278086;
Input[1470]<=14189277;
Input[1471]<=14099048;
Input[1472]<=14007410;
Input[1473]<=13914371;
Input[1474]<=13819940;
Input[1475]<=13724127;
Input[1476]<=13626942;
Input[1477]<=13528395;
Input[1478]<=13428494;
Input[1479]<=13327251;
Input[1480]<=13224675;
Input[1481]<=13120776;
Input[1482]<=13015566;
Input[1483]<=12909053;
Input[1484]<=12801250;
Input[1485]<=12692167;
Input[1486]<=12581815;
Input[1487]<=12470204;
Input[1488]<=12357347;
Input[1489]<=12243254;
Input[1490]<=12127936;
Input[1491]<=12011406;
Input[1492]<=11893674;
Input[1493]<=11774753;
Input[1494]<=11654655;
Input[1495]<=11533391;
Input[1496]<=11410974;
Input[1497]<=11287416;
Input[1498]<=11162729;
Input[1499]<=11036926;
Input[1500]<=10910019;
Input[1501]<=10782021;
Input[1502]<=10652945;
Input[1503]<=10522804;
Input[1504]<=10391610;
Input[1505]<=10259377;
Input[1506]<=10126119;
Input[1507]<=9991847;
Input[1508]<=9856577;
Input[1509]<=9720321;
Input[1510]<=9583093;
Input[1511]<=9444906;
Input[1512]<=9305775;
Input[1513]<=9165714;
Input[1514]<=9024736;
Input[1515]<=8882855;
Input[1516]<=8740087;
Input[1517]<=8596444;
Input[1518]<=8451941;
Input[1519]<=8306594;
Input[1520]<=8160415;
Input[1521]<=8013421;
Input[1522]<=7865625;
Input[1523]<=7717043;
Input[1524]<=7567689;
Input[1525]<=7417579;
Input[1526]<=7266726;
Input[1527]<=7115147;
Input[1528]<=6962857;
Input[1529]<=6809870;
Input[1530]<=6656202;
Input[1531]<=6501868;
Input[1532]<=6346885;
Input[1533]<=6191266;
Input[1534]<=6035029;
Input[1535]<=5878188;
Input[1536]<=5720759;
Input[1537]<=5562758;
Input[1538]<=5404201;
Input[1539]<=5245104;
Input[1540]<=5085482;
Input[1541]<=4925351;
Input[1542]<=4764728;
Input[1543]<=4603628;
Input[1544]<=4442068;
Input[1545]<=4280064;
Input[1546]<=4117632;
Input[1547]<=3954788;
Input[1548]<=3791549;
Input[1549]<=3627930;
Input[1550]<=3463949;
Input[1551]<=3299621;
Input[1552]<=3134964;
Input[1553]<=2969992;
Input[1554]<=2804724;
Input[1555]<=2639176;
Input[1556]<=2473363;
Input[1557]<=2307303;
Input[1558]<=2141013;
Input[1559]<=1974508;
Input[1560]<=1807806;
Input[1561]<=1640923;
Input[1562]<=1473876;
Input[1563]<=1306681;
Input[1564]<=1139356;
Input[1565]<=971917;
Input[1566]<=804381;
Input[1567]<=636764;
Input[1568]<=469084;
Input[1569]<=301357;
Input[1570]<=133600;
Input[1571]<=-34170;
Input[1572]<=-201937;
Input[1573]<=-369685;
Input[1574]<=-537395;
Input[1575]<=-705051;
Input[1576]<=-872637;
Input[1577]<=-1040136;
Input[1578]<=-1207530;
Input[1579]<=-1374804;
Input[1580]<=-1541941;
Input[1581]<=-1708923;
Input[1582]<=-1875734;
Input[1583]<=-2042358;
Input[1584]<=-2208777;
Input[1585]<=-2374976;
Input[1586]<=-2540937;
Input[1587]<=-2706644;
Input[1588]<=-2872081;
Input[1589]<=-3037230;
Input[1590]<=-3202075;
Input[1591]<=-3366600;
Input[1592]<=-3530789;
Input[1593]<=-3694624;
Input[1594]<=-3858091;
Input[1595]<=-4021171;
Input[1596]<=-4183849;
Input[1597]<=-4346109;
Input[1598]<=-4507934;
Input[1599]<=-4669308;
Input[1600]<=-4830216;
Input[1601]<=-4990640;
Input[1602]<=-5150565;
Input[1603]<=-5309976;
Input[1604]<=-5468855;
Input[1605]<=-5627187;
Input[1606]<=-5784957;
Input[1607]<=-5942148;
Input[1608]<=-6098745;
Input[1609]<=-6254733;
Input[1610]<=-6410094;
Input[1611]<=-6564815;
Input[1612]<=-6718879;
Input[1613]<=-6872271;
Input[1614]<=-7024976;
Input[1615]<=-7176979;
Input[1616]<=-7328264;
Input[1617]<=-7478816;
Input[1618]<=-7628620;
Input[1619]<=-7777662;
Input[1620]<=-7925925;
Input[1621]<=-8073396;
Input[1622]<=-8220060;
Input[1623]<=-8365902;
Input[1624]<=-8510907;
Input[1625]<=-8655061;
Input[1626]<=-8798349;
Input[1627]<=-8940758;
Input[1628]<=-9082272;
Input[1629]<=-9222879;
Input[1630]<=-9362563;
Input[1631]<=-9501311;
Input[1632]<=-9639109;
Input[1633]<=-9775942;
Input[1634]<=-9911799;
Input[1635]<=-10046664;
Input[1636]<=-10180524;
Input[1637]<=-10313367;
Input[1638]<=-10445178;
Input[1639]<=-10575944;
Input[1640]<=-10705653;
Input[1641]<=-10834292;
Input[1642]<=-10961847;
Input[1643]<=-11088305;
Input[1644]<=-11213655;
Input[1645]<=-11337884;
Input[1646]<=-11460979;
Input[1647]<=-11582928;
Input[1648]<=-11703718;
Input[1649]<=-11823338;
Input[1650]<=-11941776;
Input[1651]<=-12059020;
Input[1652]<=-12175057;
Input[1653]<=-12289878;
Input[1654]<=-12403469;
Input[1655]<=-12515820;
Input[1656]<=-12626919;
Input[1657]<=-12736756;
Input[1658]<=-12845319;
Input[1659]<=-12952597;
Input[1660]<=-13058580;
Input[1661]<=-13163258;
Input[1662]<=-13266619;
Input[1663]<=-13368653;
Input[1664]<=-13469351;
Input[1665]<=-13568702;
Input[1666]<=-13666695;
Input[1667]<=-13763322;
Input[1668]<=-13858573;
Input[1669]<=-13952438;
Input[1670]<=-14044908;
Input[1671]<=-14135973;
Input[1672]<=-14225625;
Input[1673]<=-14313854;
Input[1674]<=-14400652;
Input[1675]<=-14486009;
Input[1676]<=-14569918;
Input[1677]<=-14652371;
Input[1678]<=-14733357;
Input[1679]<=-14812871;
Input[1680]<=-14890903;
Input[1681]<=-14967447;
Input[1682]<=-15042493;
Input[1683]<=-15116035;
Input[1684]<=-15188066;
Input[1685]<=-15258578;
Input[1686]<=-15327564;
Input[1687]<=-15395017;
Input[1688]<=-15460931;
Input[1689]<=-15525299;
Input[1690]<=-15588114;
Input[1691]<=-15649370;
Input[1692]<=-15709062;
Input[1693]<=-15767182;
Input[1694]<=-15823726;
Input[1695]<=-15878688;
Input[1696]<=-15932061;
Input[1697]<=-15983842;
Input[1698]<=-16034024;
Input[1699]<=-16082602;
Input[1700]<=-16129573;
Input[1701]<=-16174930;
Input[1702]<=-16218670;
Input[1703]<=-16260789;
Input[1704]<=-16301281;
Input[1705]<=-16340143;
Input[1706]<=-16377371;
Input[1707]<=-16412961;
Input[1708]<=-16446910;
Input[1709]<=-16479214;
Input[1710]<=-16509871;
Input[1711]<=-16538876;
Input[1712]<=-16566228;
Input[1713]<=-16591923;
Input[1714]<=-16615958;
Input[1715]<=-16638333;
Input[1716]<=-16659043;
Input[1717]<=-16678087;
Input[1718]<=-16695464;
Input[1719]<=-16711171;
Input[1720]<=-16725207;
Input[1721]<=-16737571;
Input[1722]<=-16748261;
Input[1723]<=-16757276;
Input[1724]<=-16764615;
Input[1725]<=-16770278;
Input[1726]<=-16774263;
Input[1727]<=-16776572;
Input[1728]<=-16777203;
Input[1729]<=-16776156;
Input[1730]<=-16773431;
Input[1731]<=-16769029;
Input[1732]<=-16762950;
Input[1733]<=-16755195;
Input[1734]<=-16745765;
Input[1735]<=-16734660;
Input[1736]<=-16721881;
Input[1737]<=-16707430;
Input[1738]<=-16691309;
Input[1739]<=-16673518;
Input[1740]<=-16654060;
Input[1741]<=-16632937;
Input[1742]<=-16610150;
Input[1743]<=-16585703;
Input[1744]<=-16559597;
Input[1745]<=-16531835;
Input[1746]<=-16502419;
Input[1747]<=-16471354;
Input[1748]<=-16438641;
Input[1749]<=-16404285;
Input[1750]<=-16368288;
Input[1751]<=-16330654;
Input[1752]<=-16291387;
Input[1753]<=-16250491;
Input[1754]<=-16207970;
Input[1755]<=-16163829;
Input[1756]<=-16118071;
Input[1757]<=-16070701;
Input[1758]<=-16021724;
Input[1759]<=-15971145;
Input[1760]<=-15918969;
Input[1761]<=-15865201;
Input[1762]<=-15809846;
Input[1763]<=-15752910;
Input[1764]<=-15694400;
Input[1765]<=-15634319;
Input[1766]<=-15572676;
Input[1767]<=-15509475;
Input[1768]<=-15444723;
Input[1769]<=-15378427;
Input[1770]<=-15310592;
Input[1771]<=-15241227;
Input[1772]<=-15170338;
Input[1773]<=-15097932;
Input[1774]<=-15024015;
Input[1775]<=-14948597;
Input[1776]<=-14871684;
Input[1777]<=-14793283;
Input[1778]<=-14713403;
Input[1779]<=-14632052;
Input[1780]<=-14549238;
Input[1781]<=-14464969;
Input[1782]<=-14379253;
Input[1783]<=-14292099;
Input[1784]<=-14203516;
Input[1785]<=-14113513;
Input[1786]<=-14022099;
Input[1787]<=-13929282;
Input[1788]<=-13835072;
Input[1789]<=-13739479;
Input[1790]<=-13642512;
Input[1791]<=-13544181;
Input[1792]<=-13444495;
Input[1793]<=-13343465;
Input[1794]<=-13241100;
Input[1795]<=-13137412;
Input[1796]<=-13032409;
Input[1797]<=-12926104;
Input[1798]<=-12818506;
Input[1799]<=-12709626;
Input[1800]<=-12599475;
Input[1801]<=-12488064;
Input[1802]<=-12375404;
Input[1803]<=-12261507;
Input[1804]<=-12146384;
Input[1805]<=-12030046;
Input[1806]<=-11912505;
Input[1807]<=-11793772;
Input[1808]<=-11673861;
Input[1809]<=-11552782;
Input[1810]<=-11430548;
Input[1811]<=-11307170;
Input[1812]<=-11182662;
Input[1813]<=-11057036;
Input[1814]<=-10930304;
Input[1815]<=-10802479;
Input[1816]<=-10673574;
Input[1817]<=-10543602;
Input[1818]<=-10412575;
Input[1819]<=-10280507;
Input[1820]<=-10147410;
Input[1821]<=-10013299;
Input[1822]<=-9878187;
Input[1823]<=-9742087;
Input[1824]<=-9605013;
Input[1825]<=-9466978;
Input[1826]<=-9327997;
Input[1827]<=-9188083;
Input[1828]<=-9047250;
Input[1829]<=-8905512;
Input[1830]<=-8762884;
Input[1831]<=-8619379;
Input[1832]<=-8475012;
Input[1833]<=-8329798;
Input[1834]<=-8183752;
Input[1835]<=-8036886;
Input[1836]<=-7889217;
Input[1837]<=-7740759;
Input[1838]<=-7591527;
Input[1839]<=-7441536;
Input[1840]<=-7290801;
Input[1841]<=-7139336;
Input[1842]<=-6987158;
Input[1843]<=-6834281;
Input[1844]<=-6680721;
Input[1845]<=-6526492;
Input[1846]<=-6371611;
Input[1847]<=-6216093;
Input[1848]<=-6059953;
Input[1849]<=-5903207;
Input[1850]<=-5745871;
Input[1851]<=-5587960;
Input[1852]<=-5429490;
Input[1853]<=-5270478;
Input[1854]<=-5110938;
Input[1855]<=-4950888;
Input[1856]<=-4790342;
Input[1857]<=-4629317;
Input[1858]<=-4467830;
Input[1859]<=-4305895;
Input[1860]<=-4143530;
Input[1861]<=-3980751;
Input[1862]<=-3817573;
Input[1863]<=-3654014;
Input[1864]<=-3490089;
Input[1865]<=-3325816;
Input[1866]<=-3161209;
Input[1867]<=-2996287;
Input[1868]<=-2831065;
Input[1869]<=-2665560;
Input[1870]<=-2499788;
Input[1871]<=-2333767;
Input[1872]<=-2167512;
Input[1873]<=-2001040;
Input[1874]<=-1834368;
Input[1875]<=-1667513;
Input[1876]<=-1500491;
Input[1877]<=-1333319;
Input[1878]<=-1166013;
Input[1879]<=-998591;
Input[1880]<=-831070;
Input[1881]<=-663465;
Input[1882]<=-495793;
Input[1883]<=-328073;
Input[1884]<=-160319;

Signal<=0;
SigInd <=0;

end

always @( posedge control )
begin
	// Output = stored values
	
	
		Signal = Input[i];
		i=i+1;
		SigInd = !SigInd;
		if (i>SignalLength)
		begin
		i=0;
		end
end

endmodule
